* SPICE3 file created from dac.ext - technology: sky130A

X0 VN current_mirror_0/IB current_mirror_0/a_35500_32800# VN sky130_fd_pr__nfet_01v8 ad=16 pd=16 as=16 ps=12 w=4 l=12
X1 current_mirror_0/a_35500_32800# m2m_ladder_0/IOUT IOUT VN sky130_fd_pr__nfet_01v8 ad=16 pd=12 as=16 ps=16 w=4 l=12
X2 VN current_mirror_0/IB current_mirror_0/a_35500_30000# VN sky130_fd_pr__nfet_01v8 ad=16 pd=16 as=16 ps=12 w=4 l=12
X3 current_mirror_0/a_35500_30000# m2m_ladder_0/IOUT m2m_ladder_0/IOUT VN sky130_fd_pr__nfet_01v8 ad=16 pd=12 as=16 ps=16 w=4 l=12
X4 current_mirror_0/a_35500_30000# current_mirror_0/IB current_mirror_0/IB VN sky130_fd_pr__nfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X5 bias_gen_0/a_17900_29830# bias_gen_0/a_17900_29830# VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X6 VN bias_gen_0/a_15100_29900# bias_gen_0/a_17900_29830# VN sky130_fd_pr__nfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X7 bias_gen_0/a_15100_29900# bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X8 V bias_gen_0/a_15100_29900# bias_gen_0/a_15100_29900# VN sky130_fd_pr__nfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X9 V bias_gen_0/a_15100_29900# bias_gen_0/a_15100_29900# VN sky130_fd_pr__nfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X10 V bias_gen_0/a_15100_29900# bias_gen_0/a_15100_29900# VN sky130_fd_pr__nfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X11 bias_gen_0/VBP bias_gen_0/a_17900_29830# VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X12 VN bias_gen_0/a_15100_31900# bias_gen_0/a_15100_31900# VN sky130_fd_pr__nfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X13 VN bias_gen_0/a_15100_31900# bias_gen_0/VBP VN sky130_fd_pr__nfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X14 bias_gen_0/a_15100_31900# bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X15 m2m_ladder_0/a_8000_7800# m2m_ladder_0/a_5600_9530# m2m_ladder_0/IOUT VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X16 m2m_ladder_0/a_20600_7800# D2 VN VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X17 m2m_ladder_0/a_22600_9530# D1 VP VP sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X18 m2m_ladder_0/a_27000_9530# D0 VP VP sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X19 m2m_ladder_0/a_25000_13400# bias_gen_0/VBP m2m_ladder_0/a_20600_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X20 m2m_ladder_0/a_12200_7800# m2m_ladder_0/a_9800_9530# m2m_ladder_0/IOUT VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X21 m2m_ladder_0/a_3800_13400# bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X22 m2m_ladder_0/a_20600_13400# bias_gen_0/VBP m2m_ladder_0/a_16400_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X23 m2m_ladder_0/a_25000_13400# bias_gen_0/VBP m2m_ladder_0/a_20600_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X24 m2m_ladder_0/a_25000_7800# m2m_ladder_0/a_22600_9530# m2m_ladder_0/IOUT VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X25 m2m_ladder_0/a_29400_7800# m2m_ladder_0/a_27000_9530# m2m_ladder_0/IOUT VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X26 m2m_ladder_0/a_1400_9530# D6 VN VN sky130_fd_pr__nfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X27 m2m_ladder_0/a_9800_9530# D4 VP VP sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X28 m2m_ladder_0/a_3800_13400# bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X29 m2m_ladder_0/a_20600_13400# bias_gen_0/VBP m2m_ladder_0/a_16400_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X30 m2m_ladder_0/a_25000_7800# bias_gen_0/VBP m2m_ladder_0/a_20600_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X31 m2m_ladder_0/a_3800_7800# bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X32 m2m_ladder_0/a_20600_7800# bias_gen_0/VBP m2m_ladder_0/a_16400_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X33 m2m_ladder_0/a_3800_7800# D6 VN VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X34 m2m_ladder_0/a_5600_9530# D5 VN VN sky130_fd_pr__nfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X35 m2m_ladder_0/a_14000_9530# D3 VP VP sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X36 m2m_ladder_0/a_16400_13400# bias_gen_0/VBP m2m_ladder_0/a_12200_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X37 m2m_ladder_0/a_16400_13400# bias_gen_0/VBP m2m_ladder_0/a_12200_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X38 m2m_ladder_0/a_16400_7800# m2m_ladder_0/a_14000_9530# m2m_ladder_0/IOUT VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X39 m2m_ladder_0/a_8000_7800# D5 VN VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X40 m2m_ladder_0/a_22600_9530# D1 VN VN sky130_fd_pr__nfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X41 m2m_ladder_0/a_27000_9530# D0 VN VN sky130_fd_pr__nfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X42 m2m_ladder_0/a_18200_9530# D2 VP VP sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X43 m2m_ladder_0/a_16400_7800# bias_gen_0/VBP m2m_ladder_0/a_12200_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X44 m2m_ladder_0/a_29400_13400# bias_gen_0/VBP m2m_ladder_0/a_25000_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=12 as=16 ps=16 w=4 l=12
X45 m2m_ladder_0/a_12200_13400# bias_gen_0/VBP m2m_ladder_0/a_8000_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X46 m2m_ladder_0/a_29400_13400# bias_gen_0/VBP m2m_ladder_0/a_25000_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=12 as=16 ps=16 w=4 l=12
X47 m2m_ladder_0/a_20600_7800# m2m_ladder_0/a_18200_9530# m2m_ladder_0/IOUT VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X48 m2m_ladder_0/a_12200_7800# D4 VN VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X49 m2m_ladder_0/a_25000_7800# D1 VN VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X50 m2m_ladder_0/a_29400_7800# D0 VN VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X51 m2m_ladder_0/a_9800_9530# D4 VN VN sky130_fd_pr__nfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X52 m2m_ladder_0/a_12200_13400# bias_gen_0/VBP m2m_ladder_0/a_8000_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X53 m2m_ladder_0/a_29400_7800# bias_gen_0/VBP m2m_ladder_0/a_25000_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X54 m2m_ladder_0/a_12200_7800# bias_gen_0/VBP m2m_ladder_0/a_8000_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X55 m2m_ladder_0/a_1400_9530# D6 VP VP sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X56 m2m_ladder_0/a_14000_9530# D3 VN VN sky130_fd_pr__nfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X57 m2m_ladder_0/a_3800_7800# m2m_ladder_0/a_1400_9530# m2m_ladder_0/IOUT VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X58 m2m_ladder_0/a_8000_13400# bias_gen_0/VBP m2m_ladder_0/a_3800_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X59 VN bias_gen_0/VBP m2m_ladder_0/a_29400_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=12 w=4 l=12
X60 m2m_ladder_0/a_5600_9530# D5 VP VP sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X61 m2m_ladder_0/a_8000_13400# bias_gen_0/VBP m2m_ladder_0/a_3800_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X62 m2m_ladder_0/a_16400_7800# D3 VN VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X63 m2m_ladder_0/a_18200_9530# D2 VN VN sky130_fd_pr__nfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X64 VN bias_gen_0/VBP m2m_ladder_0/a_29400_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=12 w=4 l=12
X65 m2m_ladder_0/a_8000_7800# bias_gen_0/VBP m2m_ladder_0/a_3800_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X66 current_divider_0/a_27400_1800# bias_gen_0/VBP current_divider_0/a_22400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X67 current_mirror_0/IB bias_gen_0/VBP current_divider_0/a_62400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=12 w=4 l=12
X68 VN bias_gen_0/VBP current_divider_0/a_37400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X69 VP bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=993.57501 ps=1.0053k w=4 l=12
X70 VP bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X71 current_divider_0/a_17400_1800# bias_gen_0/VBP current_divider_0/a_12400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X72 VN bias_gen_0/VBP current_divider_0/a_17400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X73 VN bias_gen_0/VBP current_divider_0/a_27400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X74 VP bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X75 VN bias_gen_0/VBP current_divider_0/a_7400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X76 current_divider_0/a_7400_1800# bias_gen_0/VBP current_divider_0/a_2400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X77 current_divider_0/a_7400_1800# bias_gen_0/VBP current_divider_0/a_2400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X78 VP bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X79 VP bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X80 VP bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X81 VP bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X82 VP bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X83 VP bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X84 current_divider_0/a_62400_1800# bias_gen_0/VBP current_divider_0/a_57400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=12 as=16 ps=16 w=4 l=12
X85 VP bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X86 VP bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X87 VP bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X88 current_divider_0/a_52400_1800# bias_gen_0/VBP current_divider_0/a_47400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X89 current_divider_0/a_62400_1800# bias_gen_0/VBP current_divider_0/a_57400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=12 as=16 ps=16 w=4 l=12
X90 VP bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X91 current_divider_0/a_42400_1800# bias_gen_0/VBP current_divider_0/a_37400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X92 current_divider_0/a_52400_1800# bias_gen_0/VBP current_divider_0/a_47400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X93 VP bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X94 current_divider_0/a_22400_1800# bias_gen_0/VBP current_divider_0/a_17400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X95 current_divider_0/a_32400_1800# bias_gen_0/VBP current_divider_0/a_27400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X96 current_divider_0/a_42400_1800# bias_gen_0/VBP current_divider_0/a_37400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X97 VP bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X98 current_divider_0/a_12400_1800# bias_gen_0/VBP current_divider_0/a_7400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X99 current_divider_0/a_22400_1800# bias_gen_0/VBP current_divider_0/a_17400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X100 current_divider_0/a_32400_1800# bias_gen_0/VBP current_divider_0/a_27400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X101 current_divider_0/a_12400_1800# bias_gen_0/VBP current_divider_0/a_7400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X102 VN bias_gen_0/VBP current_divider_0/a_42400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X103 VN bias_gen_0/VBP current_divider_0/a_52400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X104 VP bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X105 VN bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X106 VN bias_gen_0/VBP current_divider_0/a_32400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X107 VN bias_gen_0/VBP current_divider_0/a_22400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X108 VN bias_gen_0/VBP current_divider_0/a_12400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X109 VP bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X110 VN bias_gen_0/VBP current_divider_0/a_2400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X111 VP bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X112 VP bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X113 VP bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X114 VP bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X115 VP bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X116 VP bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X117 current_divider_0/a_47400_1800# bias_gen_0/VBP current_divider_0/a_42400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X118 current_divider_0/a_57400_1800# bias_gen_0/VBP current_divider_0/a_52400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X119 VP bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X120 VP bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X121 current_divider_0/a_2400_1800# bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X122 current_divider_0/a_37400_1800# bias_gen_0/VBP current_divider_0/a_32400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X123 current_divider_0/a_47400_1800# bias_gen_0/VBP current_divider_0/a_42400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X124 current_divider_0/a_57400_1800# bias_gen_0/VBP current_divider_0/a_52400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X125 VP bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X126 current_divider_0/a_17400_1800# bias_gen_0/VBP current_divider_0/a_12400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X127 current_divider_0/a_27400_1800# bias_gen_0/VBP current_divider_0/a_22400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X128 current_mirror_0/IB bias_gen_0/VBP current_divider_0/a_62400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=12 w=4 l=12
X129 current_divider_0/a_2400_1800# bias_gen_0/VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X130 current_divider_0/a_37400_1800# bias_gen_0/VBP current_divider_0/a_32400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X131 VN bias_gen_0/VBP current_divider_0/a_47400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X132 VN bias_gen_0/VBP current_divider_0/a_57400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
