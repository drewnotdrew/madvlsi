* SPICE3 file created from dac.ext - technology: sky130A

.subckt current_mirror VN IB IIN IOUT
X0 VN IB a_35500_32800# VN sky130_fd_pr__nfet_01v8 ad=16 pd=16 as=16 ps=12 w=4 l=12
X1 a_35500_32800# IIN IOUT VN sky130_fd_pr__nfet_01v8 ad=16 pd=12 as=16 ps=16 w=4 l=12
X2 VN IB a_35500_30000# VN sky130_fd_pr__nfet_01v8 ad=16 pd=16 as=16 ps=12 w=4 l=12
X3 a_35500_30000# IIN IIN VN sky130_fd_pr__nfet_01v8 ad=16 pd=12 as=16 ps=16 w=4 l=12
X4 a_35500_30000# IB IB VN sky130_fd_pr__nfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
.ends

.subckt m2m_ladder VN VP D6 IIN D5 D4 D3 D2 D1 D0 VGATE IDUMP IOUT
X0 a_8000_7800# a_5600_9530# IOUT VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X1 a_20600_7800# D2 IDUMP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X2 a_22600_9530# D1 VP VP sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X3 a_27000_9530# D0 VP VP sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X4 a_25000_13400# VGATE a_20600_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X5 a_12200_7800# a_9800_9530# IOUT VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X6 a_3800_13400# VGATE IIN VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X7 a_20600_13400# VGATE a_16400_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X8 a_25000_13400# VGATE a_20600_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X9 a_25000_7800# a_22600_9530# IOUT VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X10 a_29400_7800# a_27000_9530# IOUT VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X11 a_1400_9530# D6 VN VN sky130_fd_pr__nfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X12 a_9800_9530# D4 VP VP sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X13 a_3800_13400# VGATE IIN VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X14 a_20600_13400# VGATE a_16400_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X15 a_25000_7800# VGATE a_20600_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X16 a_3800_7800# VGATE IIN VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X17 a_20600_7800# VGATE a_16400_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X18 a_3800_7800# D6 IDUMP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X19 a_5600_9530# D5 VN VN sky130_fd_pr__nfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X20 a_14000_9530# D3 VP VP sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X21 a_16400_13400# VGATE a_12200_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X22 a_16400_13400# VGATE a_12200_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X23 a_16400_7800# a_14000_9530# IOUT VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X24 a_8000_7800# D5 IDUMP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X25 a_22600_9530# D1 VN VN sky130_fd_pr__nfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X26 a_27000_9530# D0 VN VN sky130_fd_pr__nfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X27 a_18200_9530# D2 VP VP sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X28 a_16400_7800# VGATE a_12200_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X29 a_29400_13400# VGATE a_25000_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=12 as=16 ps=16 w=4 l=12
X30 a_12200_13400# VGATE a_8000_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X31 a_29400_13400# VGATE a_25000_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=12 as=16 ps=16 w=4 l=12
X32 a_20600_7800# a_18200_9530# IOUT VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X33 a_12200_7800# D4 IDUMP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X34 a_25000_7800# D1 IDUMP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X35 a_29400_7800# D0 IDUMP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X36 a_9800_9530# D4 VN VN sky130_fd_pr__nfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X37 a_12200_13400# VGATE a_8000_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X38 a_29400_7800# VGATE a_25000_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X39 a_12200_7800# VGATE a_8000_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X40 a_1400_9530# D6 VP VP sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X41 a_14000_9530# D3 VN VN sky130_fd_pr__nfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X42 a_3800_7800# a_1400_9530# IOUT VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X43 a_8000_13400# VGATE a_3800_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X44 IDUMP VGATE a_29400_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=12 w=4 l=12
X45 a_5600_9530# D5 VP VP sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X46 a_8000_13400# VGATE a_3800_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X47 a_16400_7800# D3 IDUMP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X48 a_18200_9530# D2 VN VN sky130_fd_pr__nfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X49 IDUMP VGATE a_29400_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=12 w=4 l=12
X50 a_8000_7800# VGATE a_3800_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
.ends

.subckt bias_gen VP V VN VBP
X0 a_17900_29830# a_17900_29830# VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X1 VN a_15100_29900# a_17900_29830# VN sky130_fd_pr__nfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X2 a_15100_29900# VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X3 V a_15100_29900# a_15100_29900# VN sky130_fd_pr__nfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X4 V a_15100_29900# a_15100_29900# VN sky130_fd_pr__nfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X5 V a_15100_29900# a_15100_29900# VN sky130_fd_pr__nfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X6 VBP a_17900_29830# VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X7 VN a_15100_31900# a_15100_31900# VN sky130_fd_pr__nfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X8 VN a_15100_31900# VBP VN sky130_fd_pr__nfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X9 a_15100_31900# VBP VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
.ends

.subckt current_divider VGATE VP VN IOUT
X0 a_27400_1800# VGATE a_22400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X1 IOUT VGATE a_62400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=12 w=4 l=12
X2 VN VGATE a_37400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X3 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=880 ps=880 w=4 l=12
X4 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X5 a_17400_1800# VGATE a_12400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X6 VN VGATE a_17400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X7 VN VGATE a_27400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X8 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X9 VN VGATE a_7400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X10 a_7400_1800# VGATE a_2400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X11 a_7400_1800# VGATE a_2400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X12 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X13 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X14 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X15 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X16 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X17 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X18 a_62400_1800# VGATE a_57400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=12 as=16 ps=16 w=4 l=12
X19 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X20 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X21 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X22 a_52400_1800# VGATE a_47400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X23 a_62400_1800# VGATE a_57400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=12 as=16 ps=16 w=4 l=12
X24 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X25 a_42400_1800# VGATE a_37400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X26 a_52400_1800# VGATE a_47400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X27 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X28 a_22400_1800# VGATE a_17400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X29 a_32400_1800# VGATE a_27400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X30 a_42400_1800# VGATE a_37400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X31 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X32 a_12400_1800# VGATE a_7400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X33 a_22400_1800# VGATE a_17400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X34 a_32400_1800# VGATE a_27400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X35 a_12400_1800# VGATE a_7400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X36 VN VGATE a_42400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X37 VN VGATE a_52400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X38 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X39 VN VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X40 VN VGATE a_32400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X41 VN VGATE a_22400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X42 VN VGATE a_12400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X43 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X44 VN VGATE a_2400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X45 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X46 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X47 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X48 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X49 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X50 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X51 a_47400_1800# VGATE a_42400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X52 a_57400_1800# VGATE a_52400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X53 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X54 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X55 a_2400_1800# VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X56 a_37400_1800# VGATE a_32400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X57 a_47400_1800# VGATE a_42400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X58 a_57400_1800# VGATE a_52400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X59 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X60 a_17400_1800# VGATE a_12400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X61 a_27400_1800# VGATE a_22400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X62 IOUT VGATE a_62400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=12 w=4 l=12
X63 a_2400_1800# VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X64 a_37400_1800# VGATE a_32400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X65 VN VGATE a_47400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X66 VN VGATE a_57400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
.ends

.subckt dac
Xcurrent_mirror_0 VSUBS current_mirror_0/IB current_mirror_0/IIN current_mirror_0/IOUT
+ current_mirror
Xm2m_ladder_0 VSUBS m2m_ladder_0/VP m2m_ladder_0/D6 m2m_ladder_0/IIN m2m_ladder_0/D5
+ m2m_ladder_0/D4 m2m_ladder_0/D3 m2m_ladder_0/D2 m2m_ladder_0/D1 m2m_ladder_0/D0
+ m2m_ladder_0/VGATE m2m_ladder_0/IDUMP m2m_ladder_0/IOUT m2m_ladder
Xbias_gen_0 bias_gen_0/VP bias_gen_0/V VSUBS bias_gen_0/VBP bias_gen
Xcurrent_divider_0 current_divider_0/VGATE current_divider_0/VP current_divider_0/VN
+ current_divider_0/IOUT current_divider
.ends

