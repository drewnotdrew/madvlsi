* SPICE3 file created from current_divider.ext - technology: sky130A

X0 a_27400_1800# VGATE a_22400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X1 IOUT VGATE a_62400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=12 w=4 l=12
X2 VN VGATE a_37400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X3 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=880 ps=880 w=4 l=12
X4 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X5 a_17400_1800# VGATE a_12400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X6 VN VGATE a_17400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X7 VN VGATE a_27400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X8 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X9 VN VGATE a_7400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X10 a_7400_1800# VGATE a_2400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X11 a_7400_1800# VGATE a_2400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X12 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X13 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X14 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X15 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X16 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X17 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X18 a_62400_1800# VGATE a_57400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=12 as=16 ps=16 w=4 l=12
X19 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X20 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X21 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X22 a_52400_1800# VGATE a_47400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X23 a_62400_1800# VGATE a_57400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=12 as=16 ps=16 w=4 l=12
X24 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X25 a_42400_1800# VGATE a_37400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X26 a_52400_1800# VGATE a_47400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X27 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X28 a_22400_1800# VGATE a_17400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X29 a_32400_1800# VGATE a_27400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X30 a_42400_1800# VGATE a_37400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X31 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X32 a_12400_1800# VGATE a_7400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X33 a_22400_1800# VGATE a_17400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X34 a_32400_1800# VGATE a_27400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X35 a_12400_1800# VGATE a_7400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X36 VN VGATE a_42400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X37 VN VGATE a_52400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X38 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X39 VN VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X40 VN VGATE a_32400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X41 VN VGATE a_22400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X42 VN VGATE a_12400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X43 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X44 VN VGATE a_2400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X45 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X46 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X47 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X48 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X49 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X50 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X51 a_47400_1800# VGATE a_42400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X52 a_57400_1800# VGATE a_52400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X53 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X54 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X55 a_2400_1800# VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X56 a_37400_1800# VGATE a_32400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X57 a_47400_1800# VGATE a_42400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X58 a_57400_1800# VGATE a_52400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X59 VP VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=0 ps=0 w=4 l=12
X60 a_17400_1800# VGATE a_12400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X61 a_27400_1800# VGATE a_22400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X62 IOUT VGATE a_62400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=12 w=4 l=12
X63 a_2400_1800# VGATE VP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X64 a_37400_1800# VGATE a_32400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X65 VN VGATE a_47400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X66 VN VGATE a_57400_1800# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
