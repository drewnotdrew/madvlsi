magic
tech sky130A
timestamp 1763033020
<< nmos >>
rect 16550 16400 17750 16800
rect 18550 16400 19750 16800
rect 16550 15500 17750 15900
rect 18550 15500 19750 15900
rect 16550 15000 17750 15400
<< ndiff >>
rect 16150 16700 16550 16800
rect 16150 16500 16250 16700
rect 16450 16500 16550 16700
rect 16150 16400 16550 16500
rect 17750 16700 18550 16800
rect 17750 16500 17850 16700
rect 18050 16500 18250 16700
rect 18450 16500 18550 16700
rect 17750 16400 18550 16500
rect 19750 16700 20150 16800
rect 19750 16500 19850 16700
rect 20050 16500 20150 16700
rect 19750 16400 20150 16500
rect 16150 15800 16550 15900
rect 16150 15600 16250 15800
rect 16450 15600 16550 15800
rect 16150 15500 16550 15600
rect 17750 15800 18550 15900
rect 17750 15600 17850 15800
rect 18050 15600 18250 15800
rect 18450 15600 18550 15800
rect 17750 15500 18550 15600
rect 19750 15800 20150 15900
rect 19750 15600 19850 15800
rect 20050 15600 20150 15800
rect 19750 15500 20150 15600
rect 16150 15300 16550 15400
rect 16150 15100 16250 15300
rect 16450 15100 16550 15300
rect 16150 15000 16550 15100
rect 17750 15300 18150 15400
rect 17750 15100 17850 15300
rect 18050 15100 18150 15300
rect 17750 15000 18150 15100
<< ndiffc >>
rect 16250 16500 16450 16700
rect 17850 16500 18050 16700
rect 18250 16500 18450 16700
rect 19850 16500 20050 16700
rect 16250 15600 16450 15800
rect 17850 15600 18050 15800
rect 18250 15600 18450 15800
rect 19850 15600 20050 15800
rect 16250 15100 16450 15300
rect 17850 15100 18050 15300
<< psubdiff >>
rect 16150 17150 16550 17250
rect 16150 16950 16250 17150
rect 16450 16950 16550 17150
rect 16150 16850 16550 16950
rect 17950 16250 18350 16350
rect 17950 16050 18050 16250
rect 18250 16050 18350 16250
rect 17950 15950 18350 16050
rect 19800 16250 20200 16350
rect 19800 16050 19900 16250
rect 20100 16050 20200 16250
rect 19800 15950 20200 16050
rect 16150 14400 16550 14500
rect 16150 14200 16250 14400
rect 16450 14200 16550 14400
rect 16150 14100 16550 14200
<< psubdiffcont >>
rect 16250 16950 16450 17150
rect 18050 16050 18250 16250
rect 19900 16050 20100 16250
rect 16250 14200 16450 14400
<< poly >>
rect 16550 16800 17750 16835
rect 18550 16800 19750 16835
rect 16550 16350 17750 16400
rect 16150 16250 17750 16350
rect 16150 16050 16250 16250
rect 16450 16050 17750 16250
rect 16150 15950 17750 16050
rect 16550 15900 17750 15950
rect 18550 15900 19750 16400
rect 16550 15465 17750 15500
rect 16550 15400 17750 15435
rect 16550 14950 17750 15000
rect 18550 14950 19750 15500
rect 16150 14850 19750 14950
rect 16150 14650 16250 14850
rect 16450 14650 19750 14850
rect 16150 14550 19750 14650
<< polycont >>
rect 16250 16050 16450 16250
rect 16250 14650 16450 14850
<< locali >>
rect 16150 17150 20200 17250
rect 16150 16950 16250 17150
rect 16450 16950 20200 17150
rect 16150 16850 20200 16950
rect 19800 16800 20200 16850
rect 16150 16700 16550 16800
rect 16150 16500 16250 16700
rect 16450 16500 16550 16700
rect 16150 16400 16550 16500
rect 17750 16700 18550 16800
rect 17750 16500 17850 16700
rect 18050 16500 18250 16700
rect 18450 16500 18550 16700
rect 17750 16400 18550 16500
rect 19750 16700 20200 16800
rect 19750 16500 19850 16700
rect 20050 16500 20200 16700
rect 19750 16400 20200 16500
rect 19800 16350 20200 16400
rect 16150 16250 16550 16350
rect 16150 16050 16250 16250
rect 16450 16050 16550 16250
rect 16150 15800 16550 16050
rect 17950 16250 20200 16350
rect 17950 16050 18050 16250
rect 18250 16050 19900 16250
rect 20100 16050 20200 16250
rect 17950 15950 20200 16050
rect 19800 15900 20200 15950
rect 16150 15600 16250 15800
rect 16450 15600 16550 15800
rect 16150 15500 16550 15600
rect 17750 15800 18550 15900
rect 17750 15600 17850 15800
rect 18050 15600 18250 15800
rect 18450 15600 18550 15800
rect 17750 15500 18550 15600
rect 19750 15800 20200 15900
rect 19750 15600 19850 15800
rect 20050 15600 20200 15800
rect 19750 15500 20200 15600
rect 17950 15400 18350 15500
rect 16150 15300 16550 15400
rect 16150 15100 16250 15300
rect 16450 15100 16550 15300
rect 16150 14850 16550 15100
rect 17750 15300 18350 15400
rect 17750 15100 17850 15300
rect 18050 15100 18350 15300
rect 17750 15000 18350 15100
rect 16150 14650 16250 14850
rect 16450 14650 16550 14850
rect 16150 14550 16550 14650
rect 19800 14500 20200 15500
rect 16150 14400 20200 14500
rect 16150 14200 16250 14400
rect 16450 14200 20200 14400
rect 16150 14100 20200 14200
<< labels >>
rlabel locali 20200 14100 20200 17250 3 VN
port 1 e
rlabel locali 16150 14550 16150 15400 7 IB
port 2 w
rlabel locali 16150 15500 16150 16350 7 IIN
port 3 w
rlabel locali 16150 16400 16150 16800 7 IOUT
port 4 w
<< end >>
