magic
tech sky130A
timestamp 1760007314
<< nwell >>
rect 380 490 860 730
rect 380 470 565 490
rect 380 180 525 470
<< nmos >>
rect 650 405 665 455
rect 650 265 665 315
rect 485 -55 500 145
rect 555 95 570 145
rect 555 -55 570 -5
rect 700 115 715 165
rect 700 -40 715 10
<< pmos >>
rect 445 645 460 695
rect 445 490 460 540
rect 445 340 460 390
rect 445 200 460 250
rect 690 510 705 710
rect 760 660 775 710
rect 760 510 775 560
<< ndiff >>
rect 605 440 650 455
rect 605 420 615 440
rect 635 420 650 440
rect 605 405 650 420
rect 665 440 710 455
rect 665 420 680 440
rect 700 420 710 440
rect 665 405 710 420
rect 605 300 650 315
rect 605 280 615 300
rect 635 280 650 300
rect 605 265 650 280
rect 665 300 710 315
rect 665 280 680 300
rect 700 280 710 300
rect 665 265 710 280
rect 440 135 485 145
rect 440 -45 450 135
rect 470 -45 485 135
rect 440 -55 485 -45
rect 500 135 555 145
rect 500 -45 515 135
rect 535 95 555 135
rect 570 130 615 145
rect 570 110 585 130
rect 605 110 615 130
rect 570 95 615 110
rect 535 -5 545 95
rect 535 -45 555 -5
rect 500 -55 555 -45
rect 570 -20 615 -5
rect 570 -40 585 -20
rect 605 -40 615 -20
rect 570 -55 615 -40
rect 655 150 700 165
rect 655 130 665 150
rect 685 130 700 150
rect 655 115 700 130
rect 715 150 760 165
rect 715 130 730 150
rect 750 130 760 150
rect 715 115 760 130
rect 655 -5 700 10
rect 655 -25 665 -5
rect 685 -25 700 -5
rect 655 -40 700 -25
rect 715 -5 760 10
rect 715 -25 730 -5
rect 750 -25 760 -5
rect 715 -40 760 -25
<< pdiff >>
rect 645 700 690 710
rect 400 680 445 695
rect 400 660 410 680
rect 430 660 445 680
rect 400 645 445 660
rect 460 680 505 695
rect 460 660 475 680
rect 495 660 505 680
rect 460 645 505 660
rect 400 525 445 540
rect 400 505 410 525
rect 430 505 445 525
rect 400 490 445 505
rect 460 525 505 540
rect 460 505 475 525
rect 495 505 505 525
rect 460 490 505 505
rect 400 375 445 390
rect 400 355 410 375
rect 430 355 445 375
rect 400 340 445 355
rect 460 375 505 390
rect 460 355 475 375
rect 495 355 505 375
rect 460 340 505 355
rect 400 235 445 250
rect 400 215 410 235
rect 430 215 445 235
rect 400 200 445 215
rect 460 235 505 250
rect 460 215 475 235
rect 495 215 505 235
rect 460 200 505 215
rect 645 515 655 700
rect 675 515 690 700
rect 645 510 690 515
rect 705 700 760 710
rect 705 515 720 700
rect 740 660 760 700
rect 775 695 820 710
rect 775 675 790 695
rect 810 675 820 695
rect 775 660 820 675
rect 740 560 750 660
rect 740 515 760 560
rect 705 510 760 515
rect 775 545 820 560
rect 775 525 790 545
rect 810 525 820 545
rect 775 510 820 525
<< ndiffc >>
rect 615 420 635 440
rect 680 420 700 440
rect 615 280 635 300
rect 680 280 700 300
rect 450 -45 470 135
rect 515 -45 535 135
rect 585 110 605 130
rect 585 -40 605 -20
rect 665 130 685 150
rect 730 130 750 150
rect 665 -25 685 -5
rect 730 -25 750 -5
<< pdiffc >>
rect 410 660 430 680
rect 475 660 495 680
rect 410 505 430 525
rect 475 505 495 525
rect 410 355 430 375
rect 475 355 495 375
rect 410 215 430 235
rect 475 215 495 235
rect 655 515 675 700
rect 720 515 740 700
rect 790 675 810 695
rect 790 525 810 545
<< psubdiff >>
rect 760 150 800 165
rect 760 130 770 150
rect 790 130 800 150
rect 760 115 800 130
<< nsubdiff >>
rect 605 695 645 710
rect 505 525 545 540
rect 505 505 515 525
rect 535 505 545 525
rect 505 490 545 505
rect 605 525 615 695
rect 635 525 645 695
rect 605 510 645 525
<< psubdiffcont >>
rect 770 130 790 150
<< nsubdiffcont >>
rect 515 505 535 525
rect 615 525 635 695
<< poly >>
rect 690 710 705 725
rect 760 720 850 735
rect 760 710 775 720
rect 445 695 460 710
rect 445 625 460 645
rect 420 615 460 625
rect 420 595 430 615
rect 450 600 460 615
rect 450 595 580 600
rect 420 585 580 595
rect 445 540 460 560
rect 445 470 460 490
rect 445 460 485 470
rect 445 440 455 460
rect 475 445 485 460
rect 475 440 540 445
rect 445 430 540 440
rect 445 390 460 405
rect 445 315 460 340
rect 420 305 460 315
rect 420 285 430 305
rect 450 285 460 305
rect 420 275 460 285
rect 445 250 460 275
rect 445 180 460 200
rect 445 165 500 180
rect 485 145 500 165
rect 525 170 540 430
rect 565 235 580 585
rect 760 645 775 660
rect 760 610 810 620
rect 760 590 780 610
rect 800 590 810 610
rect 760 580 810 590
rect 760 560 775 580
rect 690 490 705 510
rect 760 500 775 510
rect 650 475 705 490
rect 730 485 775 500
rect 650 455 665 475
rect 650 380 665 405
rect 625 370 665 380
rect 625 350 635 370
rect 655 350 665 370
rect 625 340 665 350
rect 650 315 665 340
rect 650 250 665 265
rect 730 240 745 485
rect 835 455 850 720
rect 565 225 605 235
rect 565 205 575 225
rect 595 215 605 225
rect 690 230 745 240
rect 595 205 645 215
rect 565 200 645 205
rect 690 210 700 230
rect 720 210 745 230
rect 770 445 850 455
rect 770 425 780 445
rect 800 440 850 445
rect 800 425 810 440
rect 770 415 810 425
rect 690 200 730 210
rect 565 195 605 200
rect 525 155 570 170
rect 555 145 570 155
rect 555 75 570 95
rect 555 65 605 75
rect 555 45 575 65
rect 595 45 605 65
rect 555 35 605 45
rect 555 -5 570 10
rect 485 -70 500 -55
rect 555 -65 570 -55
rect 630 -65 645 200
rect 700 165 715 200
rect 770 195 785 415
rect 770 180 835 195
rect 700 95 715 115
rect 820 70 835 180
rect 675 60 835 70
rect 675 40 685 60
rect 705 55 835 60
rect 705 40 715 55
rect 675 30 715 40
rect 700 10 715 30
rect 700 -55 715 -40
rect 555 -80 645 -65
<< polycont >>
rect 430 595 450 615
rect 455 440 475 460
rect 430 285 450 305
rect 780 590 800 610
rect 635 350 655 370
rect 575 205 595 225
rect 700 210 720 230
rect 780 425 800 445
rect 575 45 595 65
rect 685 40 705 60
<< locali >>
rect 420 715 545 735
rect 420 695 440 715
rect 400 680 440 695
rect 400 660 410 680
rect 430 660 440 680
rect 400 645 440 660
rect 465 680 505 695
rect 465 660 475 680
rect 495 660 505 680
rect 465 645 505 660
rect 420 615 460 625
rect 420 595 430 615
rect 450 595 460 615
rect 420 585 460 595
rect 420 540 440 585
rect 485 540 505 645
rect 525 605 545 715
rect 605 700 685 710
rect 605 695 655 700
rect 525 585 585 605
rect 400 525 440 540
rect 400 505 410 525
rect 430 505 440 525
rect 400 490 440 505
rect 465 525 545 540
rect 465 505 475 525
rect 495 505 515 525
rect 535 505 545 525
rect 465 490 545 505
rect 445 460 485 470
rect 400 390 420 455
rect 445 440 455 460
rect 475 455 485 460
rect 565 455 585 585
rect 605 525 615 695
rect 635 525 655 695
rect 605 515 655 525
rect 675 515 685 700
rect 605 510 685 515
rect 710 700 750 710
rect 710 515 720 700
rect 740 515 750 700
rect 780 695 820 710
rect 780 675 790 695
rect 810 675 820 695
rect 780 660 820 675
rect 790 620 810 660
rect 770 610 810 620
rect 770 590 780 610
rect 800 590 810 610
rect 770 580 810 590
rect 710 510 750 515
rect 780 545 820 560
rect 780 525 790 545
rect 810 525 820 545
rect 780 510 820 525
rect 780 455 800 510
rect 475 440 645 455
rect 445 435 615 440
rect 445 430 485 435
rect 465 390 485 430
rect 605 420 615 435
rect 635 420 645 440
rect 605 405 645 420
rect 670 445 860 455
rect 670 440 780 445
rect 670 420 680 440
rect 700 435 780 440
rect 700 420 710 435
rect 670 405 710 420
rect 770 425 780 435
rect 800 435 860 445
rect 800 425 810 435
rect 770 415 810 425
rect 400 375 440 390
rect 400 355 410 375
rect 430 355 440 375
rect 400 340 440 355
rect 465 375 505 390
rect 465 355 475 375
rect 495 355 505 375
rect 465 340 505 355
rect 545 370 830 380
rect 545 360 635 370
rect 420 305 460 315
rect 400 285 430 305
rect 450 295 460 305
rect 545 295 565 360
rect 625 350 635 360
rect 655 360 830 370
rect 655 350 665 360
rect 625 340 665 350
rect 450 285 565 295
rect 420 275 565 285
rect 605 300 645 315
rect 605 280 615 300
rect 635 280 645 300
rect 605 265 645 280
rect 670 300 790 315
rect 670 280 680 300
rect 700 295 790 300
rect 700 280 710 295
rect 670 265 710 280
rect 400 235 440 250
rect 400 215 410 235
rect 430 215 440 235
rect 400 200 440 215
rect 465 235 505 250
rect 605 235 625 265
rect 465 215 475 235
rect 495 220 505 235
rect 565 225 625 235
rect 565 220 575 225
rect 495 215 575 220
rect 465 205 575 215
rect 595 215 625 225
rect 690 240 710 265
rect 690 230 730 240
rect 595 205 605 215
rect 465 200 605 205
rect 690 210 700 230
rect 720 210 730 230
rect 690 200 730 210
rect 770 220 790 295
rect 810 305 830 360
rect 810 285 860 305
rect 770 200 860 220
rect 565 195 605 200
rect 585 145 605 195
rect 655 150 695 165
rect 400 135 480 145
rect 400 130 450 135
rect 400 -40 410 130
rect 430 -40 450 130
rect 400 -45 450 -40
rect 470 -45 480 135
rect 400 -55 480 -45
rect 505 135 545 145
rect 505 -45 515 135
rect 535 -45 545 135
rect 575 130 615 145
rect 575 110 585 130
rect 605 110 615 130
rect 655 130 665 150
rect 685 130 695 150
rect 655 115 695 130
rect 720 150 800 165
rect 720 130 730 150
rect 750 130 770 150
rect 790 130 800 150
rect 720 115 800 130
rect 575 95 615 110
rect 565 65 605 75
rect 565 45 575 65
rect 595 45 605 65
rect 565 35 605 45
rect 585 -5 605 35
rect 675 70 695 115
rect 675 60 715 70
rect 675 40 685 60
rect 705 40 715 60
rect 675 30 715 40
rect 740 10 760 115
rect 820 70 840 200
rect 655 -5 695 10
rect 505 -55 545 -45
rect 575 -20 615 -5
rect 575 -40 585 -20
rect 605 -40 615 -20
rect 655 -25 665 -5
rect 685 -25 695 -5
rect 655 -40 695 -25
rect 720 -5 760 10
rect 720 -25 730 -5
rect 750 -25 760 -5
rect 720 -40 760 -25
rect 780 50 840 70
rect 575 -55 615 -40
rect 675 -60 695 -40
rect 780 -60 800 50
rect 675 -80 800 -60
<< viali >>
rect 515 505 535 525
rect 615 525 635 695
rect 410 -40 430 130
rect 770 130 790 150
<< metal1 >>
rect 400 695 860 735
rect 400 525 615 695
rect 635 525 860 695
rect 400 505 515 525
rect 535 505 860 525
rect 400 490 860 505
rect 400 150 860 165
rect 400 130 770 150
rect 790 130 860 150
rect 400 -40 410 130
rect 430 -40 860 130
rect 400 -80 860 -40
<< labels >>
rlabel locali 400 285 400 305 7 clk
port 2 w
rlabel locali 400 200 400 220 7 Dn
port 7 w
rlabel locali 400 435 400 455 7 D
port 6 w
rlabel locali 860 200 860 220 3 Qn
port 5 e
rlabel locali 860 435 860 455 3 Q
port 4 e
rlabel metal1 400 -80 400 -60 7 VN
port 3 w
rlabel metal1 400 715 400 735 7 VP
port 1 w
<< end >>
