magic
tech sky130A
timestamp 1760277467
<< nwell >>
rect 70 490 570 730
rect 305 470 530 490
rect 305 180 450 470
<< nmos >>
rect 155 405 170 455
rect 155 265 170 315
rect 155 115 170 165
rect 155 -40 170 10
rect 400 -55 415 145
rect 470 95 485 145
rect 470 -55 485 -5
<< pmos >>
rect 195 510 210 710
rect 265 660 280 710
rect 265 510 280 560
rect 410 645 425 695
rect 410 490 425 540
rect 370 340 385 390
rect 370 200 385 250
<< ndiff >>
rect 110 440 155 455
rect 110 420 120 440
rect 140 420 155 440
rect 110 405 155 420
rect 170 440 215 455
rect 170 420 185 440
rect 205 420 215 440
rect 170 405 215 420
rect 110 300 155 315
rect 110 280 120 300
rect 140 280 155 300
rect 110 265 155 280
rect 170 300 215 315
rect 170 280 185 300
rect 205 280 215 300
rect 170 265 215 280
rect 110 150 155 165
rect 110 130 120 150
rect 140 130 155 150
rect 110 115 155 130
rect 170 150 215 165
rect 170 130 185 150
rect 205 130 215 150
rect 170 115 215 130
rect 355 135 400 145
rect 110 -5 155 10
rect 110 -25 120 -5
rect 140 -25 155 -5
rect 110 -40 155 -25
rect 170 -5 215 10
rect 170 -25 185 -5
rect 205 -25 215 -5
rect 170 -40 215 -25
rect 355 -45 365 135
rect 385 -45 400 135
rect 355 -55 400 -45
rect 415 135 470 145
rect 415 -45 430 135
rect 450 95 470 135
rect 485 130 530 145
rect 485 110 500 130
rect 520 110 530 130
rect 485 95 530 110
rect 450 -5 460 95
rect 450 -45 470 -5
rect 415 -55 470 -45
rect 485 -20 530 -5
rect 485 -40 500 -20
rect 520 -40 530 -20
rect 485 -55 530 -40
<< pdiff >>
rect 150 700 195 710
rect 150 515 160 700
rect 180 515 195 700
rect 150 510 195 515
rect 210 700 265 710
rect 210 515 225 700
rect 245 660 265 700
rect 280 695 325 710
rect 280 675 295 695
rect 315 675 325 695
rect 280 660 325 675
rect 245 560 255 660
rect 245 515 265 560
rect 210 510 265 515
rect 280 545 325 560
rect 280 525 295 545
rect 315 525 325 545
rect 280 510 325 525
rect 365 680 410 695
rect 365 660 375 680
rect 395 660 410 680
rect 365 645 410 660
rect 425 680 470 695
rect 425 660 440 680
rect 460 660 470 680
rect 425 645 470 660
rect 365 525 410 540
rect 365 505 375 525
rect 395 505 410 525
rect 365 490 410 505
rect 425 525 470 540
rect 425 505 440 525
rect 460 505 470 525
rect 425 490 470 505
rect 325 375 370 390
rect 325 355 335 375
rect 355 355 370 375
rect 325 340 370 355
rect 385 375 430 390
rect 385 355 400 375
rect 420 355 430 375
rect 385 340 430 355
rect 325 235 370 250
rect 325 215 335 235
rect 355 215 370 235
rect 325 200 370 215
rect 385 235 430 250
rect 385 215 400 235
rect 420 215 430 235
rect 385 200 430 215
<< ndiffc >>
rect 120 420 140 440
rect 185 420 205 440
rect 120 280 140 300
rect 185 280 205 300
rect 120 130 140 150
rect 185 130 205 150
rect 120 -25 140 -5
rect 185 -25 205 -5
rect 365 -45 385 135
rect 430 -45 450 135
rect 500 110 520 130
rect 500 -40 520 -20
<< pdiffc >>
rect 160 515 180 700
rect 225 515 245 700
rect 295 675 315 695
rect 295 525 315 545
rect 375 660 395 680
rect 440 660 460 680
rect 375 505 395 525
rect 440 505 460 525
rect 335 355 355 375
rect 400 355 420 375
rect 335 215 355 235
rect 400 215 420 235
<< psubdiff >>
rect 215 150 255 165
rect 215 130 225 150
rect 245 130 255 150
rect 215 115 255 130
<< nsubdiff >>
rect 110 695 150 710
rect 110 525 120 695
rect 140 525 150 695
rect 110 510 150 525
rect 470 525 510 540
rect 470 505 480 525
rect 500 505 510 525
rect 470 490 510 505
<< psubdiffcont >>
rect 225 130 245 150
<< nsubdiffcont >>
rect 120 525 140 695
rect 480 505 500 525
<< poly >>
rect 195 710 210 725
rect 265 720 355 735
rect 265 710 280 720
rect 265 645 280 660
rect 265 610 315 620
rect 265 590 285 610
rect 305 590 315 610
rect 265 580 315 590
rect 265 560 280 580
rect 195 490 210 510
rect 265 500 280 510
rect 340 500 355 720
rect 410 695 425 710
rect 410 625 425 645
rect 385 615 425 625
rect 385 595 395 615
rect 415 600 425 615
rect 415 595 545 600
rect 385 585 545 595
rect 410 540 425 560
rect 155 475 210 490
rect 235 485 280 500
rect 315 485 355 500
rect 155 455 170 475
rect 155 380 170 405
rect 130 370 170 380
rect 130 350 140 370
rect 160 350 170 370
rect 130 340 170 350
rect 155 315 170 340
rect 155 250 170 265
rect 235 240 250 485
rect 315 455 330 485
rect 410 470 425 490
rect 530 470 545 585
rect 195 230 250 240
rect 195 215 205 230
rect 155 210 205 215
rect 225 210 250 230
rect 275 445 330 455
rect 275 425 285 445
rect 305 425 330 445
rect 370 460 425 470
rect 370 440 380 460
rect 400 445 425 460
rect 490 455 545 470
rect 400 440 465 445
rect 370 430 465 440
rect 275 415 330 425
rect 155 200 235 210
rect 155 165 170 200
rect 155 100 170 115
rect 275 70 290 415
rect 370 390 385 405
rect 370 315 385 340
rect 345 305 385 315
rect 345 285 355 305
rect 375 285 385 305
rect 345 275 385 285
rect 370 250 385 275
rect 370 180 385 200
rect 450 180 465 430
rect 490 235 505 455
rect 490 225 550 235
rect 490 220 520 225
rect 510 205 520 220
rect 540 210 550 225
rect 540 205 560 210
rect 510 195 560 205
rect 370 165 415 180
rect 450 165 485 180
rect 400 145 415 165
rect 470 145 485 165
rect 130 60 290 70
rect 130 40 140 60
rect 160 55 290 60
rect 160 40 170 55
rect 130 30 170 40
rect 155 10 170 30
rect 155 -55 170 -40
rect 470 75 485 95
rect 470 65 520 75
rect 470 45 490 65
rect 510 45 520 65
rect 470 35 520 45
rect 470 -5 485 10
rect 400 -70 415 -55
rect 470 -65 485 -55
rect 545 -65 560 195
rect 470 -80 560 -65
<< polycont >>
rect 285 590 305 610
rect 395 595 415 615
rect 140 350 160 370
rect 205 210 225 230
rect 285 425 305 445
rect 380 440 400 460
rect 355 285 375 305
rect 520 205 540 225
rect 140 40 160 60
rect 490 45 510 65
<< locali >>
rect 385 715 510 735
rect 110 700 190 710
rect 110 695 160 700
rect 110 525 120 695
rect 140 525 160 695
rect 110 515 160 525
rect 180 515 190 700
rect 110 510 190 515
rect 215 700 255 710
rect 215 515 225 700
rect 245 515 255 700
rect 285 695 325 710
rect 385 695 405 715
rect 285 675 295 695
rect 315 675 325 695
rect 285 660 325 675
rect 365 680 405 695
rect 365 660 375 680
rect 395 660 405 680
rect 295 620 315 660
rect 365 645 405 660
rect 430 680 470 695
rect 430 660 440 680
rect 460 660 470 680
rect 430 645 470 660
rect 275 610 315 620
rect 275 590 285 610
rect 305 590 315 610
rect 275 580 315 590
rect 385 615 425 625
rect 385 595 395 615
rect 415 595 425 615
rect 385 585 425 595
rect 215 510 255 515
rect 285 545 325 560
rect 285 525 295 545
rect 315 525 325 545
rect 385 540 405 585
rect 450 540 470 645
rect 490 605 510 715
rect 490 585 550 605
rect 285 510 325 525
rect 365 525 405 540
rect 285 455 305 510
rect 365 505 375 525
rect 395 505 405 525
rect 365 490 405 505
rect 430 525 510 540
rect 430 505 440 525
rect 460 505 480 525
rect 500 505 510 525
rect 430 490 510 505
rect 370 460 410 470
rect 70 440 150 455
rect 70 435 120 440
rect 110 420 120 435
rect 140 420 150 440
rect 110 405 150 420
rect 175 445 315 455
rect 175 440 285 445
rect 175 420 185 440
rect 205 435 285 440
rect 205 420 215 435
rect 175 405 215 420
rect 275 425 285 435
rect 305 435 315 445
rect 370 440 380 460
rect 400 455 410 460
rect 530 455 550 585
rect 400 440 570 455
rect 370 435 570 440
rect 305 425 345 435
rect 370 430 410 435
rect 275 415 345 425
rect 325 390 345 415
rect 390 390 410 430
rect 70 370 275 380
rect 70 360 140 370
rect 130 350 140 360
rect 160 360 275 370
rect 160 350 170 360
rect 130 340 170 350
rect 255 325 275 360
rect 325 375 365 390
rect 325 355 335 375
rect 355 355 365 375
rect 325 340 365 355
rect 390 375 430 390
rect 390 355 400 375
rect 420 355 430 375
rect 390 340 430 355
rect 470 360 570 380
rect 110 300 150 315
rect 110 285 120 300
rect 70 280 120 285
rect 140 280 150 300
rect 70 265 150 280
rect 175 300 215 315
rect 255 305 315 325
rect 345 305 385 315
rect 175 280 185 300
rect 205 285 215 300
rect 295 285 355 305
rect 375 295 385 305
rect 470 295 490 360
rect 375 285 490 295
rect 205 280 275 285
rect 175 265 275 280
rect 345 275 490 285
rect 70 235 90 265
rect 195 240 215 265
rect 195 230 235 240
rect 195 210 205 230
rect 225 210 235 230
rect 195 200 235 210
rect 255 205 275 265
rect 530 265 570 285
rect 325 235 365 250
rect 325 215 335 235
rect 355 215 365 235
rect 255 185 295 205
rect 325 200 365 215
rect 390 235 430 250
rect 530 235 550 265
rect 390 215 400 235
rect 420 220 430 235
rect 510 225 550 235
rect 510 220 520 225
rect 420 215 520 220
rect 390 205 520 215
rect 540 205 550 225
rect 390 200 550 205
rect 110 150 150 165
rect 110 130 120 150
rect 140 130 150 150
rect 110 115 150 130
rect 175 150 255 165
rect 175 130 185 150
rect 205 130 225 150
rect 245 130 255 150
rect 175 115 255 130
rect 130 70 150 115
rect 130 60 170 70
rect 130 40 140 60
rect 160 40 170 60
rect 130 30 170 40
rect 195 10 215 115
rect 275 70 295 185
rect 510 195 550 200
rect 510 145 530 195
rect 110 -5 150 10
rect 110 -25 120 -5
rect 140 -25 150 -5
rect 110 -40 150 -25
rect 175 -5 215 10
rect 175 -25 185 -5
rect 205 -25 215 -5
rect 175 -40 215 -25
rect 235 50 295 70
rect 315 135 395 145
rect 315 130 365 135
rect 130 -60 150 -40
rect 235 -60 255 50
rect 315 -40 325 130
rect 345 -40 365 130
rect 315 -45 365 -40
rect 385 -45 395 135
rect 315 -55 395 -45
rect 420 135 460 145
rect 420 -45 430 135
rect 450 -45 460 135
rect 490 130 530 145
rect 490 110 500 130
rect 520 110 530 130
rect 490 95 530 110
rect 480 65 520 75
rect 480 45 490 65
rect 510 45 520 65
rect 480 35 520 45
rect 500 -5 520 35
rect 420 -55 460 -45
rect 490 -20 530 -5
rect 490 -40 500 -20
rect 520 -40 530 -20
rect 490 -55 530 -40
rect 130 -80 255 -60
<< viali >>
rect 120 525 140 695
rect 480 505 500 525
rect 225 130 245 150
rect 325 -40 345 130
<< metal1 >>
rect 70 695 570 735
rect 70 525 120 695
rect 140 525 570 695
rect 70 505 480 525
rect 500 505 570 525
rect 70 490 570 505
rect 70 150 560 165
rect 70 130 225 150
rect 245 130 560 150
rect 70 -40 325 130
rect 345 -40 560 130
rect 70 -80 560 -40
<< labels >>
rlabel metal1 70 715 70 735 7 VP
port 1 w
rlabel locali 70 435 70 455 7 D
port 2 w
rlabel locali 70 360 70 380 7 clk
port 3 w
rlabel locali 70 235 70 255 7 Dn
port 4 w
rlabel metal1 70 -80 70 -60 7 VN
port 5 w
rlabel locali 570 265 570 285 3 Qn
port 6 e
rlabel locali 570 435 570 455 3 Q
port 7 e
<< end >>
