magic
tech sky130A
timestamp 1759973783
<< error_p >>
rect 690 557 710 560
rect 515 522 535 525
rect 515 508 518 522
rect 532 508 535 522
rect 515 505 535 508
rect 690 393 693 557
rect 707 393 710 557
rect 690 390 710 393
rect 410 127 430 130
rect 410 -37 413 127
rect 427 -37 430 127
rect 795 12 815 15
rect 795 -2 798 12
rect 812 -2 815 12
rect 795 -5 815 -2
rect 410 -40 430 -37
<< nwell >>
rect 650 560 920 595
rect 380 470 920 560
rect 380 180 525 470
rect 655 360 920 470
rect 660 355 920 360
<< nmos >>
rect 725 270 740 320
rect 485 -55 500 145
rect 555 95 570 145
rect 555 -55 570 -5
rect 725 130 740 180
rect 725 -20 740 30
rect 870 -20 885 30
<< pmos >>
rect 445 490 460 540
rect 590 490 605 540
rect 445 340 460 390
rect 445 200 460 250
rect 765 375 780 575
rect 835 525 850 575
rect 835 375 850 425
<< ndiff >>
rect 680 305 725 320
rect 680 285 690 305
rect 710 285 725 305
rect 680 270 725 285
rect 740 305 785 320
rect 740 285 755 305
rect 775 285 785 305
rect 740 270 785 285
rect 440 135 485 145
rect 440 -45 450 135
rect 470 -45 485 135
rect 440 -55 485 -45
rect 500 135 555 145
rect 500 -45 515 135
rect 535 95 555 135
rect 570 130 615 145
rect 570 110 585 130
rect 605 110 615 130
rect 570 95 615 110
rect 535 -5 545 95
rect 535 -45 555 -5
rect 500 -55 555 -45
rect 570 -20 615 -5
rect 570 -40 585 -20
rect 605 -40 615 -20
rect 570 -55 615 -40
rect 680 165 725 180
rect 680 145 690 165
rect 710 145 725 165
rect 680 130 725 145
rect 740 165 785 180
rect 740 145 755 165
rect 775 145 785 165
rect 740 130 785 145
rect 680 15 725 30
rect 680 -5 690 15
rect 710 -5 725 15
rect 680 -20 725 -5
rect 740 15 785 30
rect 825 15 870 30
rect 740 -5 755 15
rect 775 -5 785 15
rect 825 -5 835 15
rect 855 -5 870 15
rect 740 -20 785 -5
rect 825 -20 870 -5
rect 885 15 930 30
rect 885 -5 900 15
rect 920 -5 930 15
rect 885 -20 930 -5
<< pdiff >>
rect 720 565 765 575
rect 400 525 445 540
rect 400 505 410 525
rect 430 505 445 525
rect 400 490 445 505
rect 460 525 505 540
rect 545 525 590 540
rect 460 505 475 525
rect 495 505 505 525
rect 545 505 555 525
rect 575 505 590 525
rect 460 490 505 505
rect 545 490 590 505
rect 605 525 650 540
rect 605 505 620 525
rect 640 505 650 525
rect 605 490 650 505
rect 400 375 445 390
rect 400 355 410 375
rect 430 355 445 375
rect 400 340 445 355
rect 460 375 505 390
rect 460 355 475 375
rect 495 355 505 375
rect 460 340 505 355
rect 400 235 445 250
rect 400 215 410 235
rect 430 215 445 235
rect 400 200 445 215
rect 460 235 505 250
rect 460 215 475 235
rect 495 215 505 235
rect 460 200 505 215
rect 720 380 730 565
rect 750 380 765 565
rect 720 375 765 380
rect 780 565 835 575
rect 780 380 795 565
rect 815 525 835 565
rect 850 560 895 575
rect 850 540 865 560
rect 885 540 895 560
rect 850 525 895 540
rect 815 425 825 525
rect 815 380 835 425
rect 780 375 835 380
rect 850 410 895 425
rect 850 390 865 410
rect 885 390 895 410
rect 850 375 895 390
<< ndiffc >>
rect 690 285 710 305
rect 755 285 775 305
rect 450 -45 470 135
rect 515 -45 535 135
rect 585 110 605 130
rect 585 -40 605 -20
rect 690 145 710 165
rect 755 145 775 165
rect 690 -5 710 15
rect 755 -5 775 15
rect 835 -5 855 15
rect 900 -5 920 15
<< pdiffc >>
rect 410 505 430 525
rect 475 505 495 525
rect 555 505 575 525
rect 620 505 640 525
rect 410 355 430 375
rect 475 355 495 375
rect 410 215 430 235
rect 475 215 495 235
rect 730 380 750 565
rect 795 380 815 565
rect 865 540 885 560
rect 865 390 885 410
<< psubdiff >>
rect 785 15 825 30
rect 785 -5 795 15
rect 815 -5 825 15
rect 785 -20 825 -5
<< nsubdiff >>
rect 680 560 720 575
rect 505 525 545 540
rect 505 505 515 525
rect 535 505 545 525
rect 505 490 545 505
rect 680 390 690 560
rect 710 390 720 560
rect 680 375 720 390
<< psubdiffcont >>
rect 795 -5 815 15
<< nsubdiffcont >>
rect 515 505 535 525
rect 690 390 710 560
<< poly >>
rect 565 590 605 600
rect 565 570 575 590
rect 595 570 605 590
rect 765 575 780 590
rect 835 585 925 600
rect 835 575 850 585
rect 565 560 605 570
rect 445 540 460 555
rect 590 540 605 560
rect 445 470 460 490
rect 590 480 605 490
rect 445 460 485 470
rect 445 440 455 460
rect 475 445 485 460
rect 565 465 605 480
rect 475 440 540 445
rect 445 430 540 440
rect 445 390 460 405
rect 445 315 460 340
rect 420 305 460 315
rect 420 285 430 305
rect 450 285 460 305
rect 420 275 460 285
rect 445 250 460 275
rect 445 180 460 200
rect 445 165 500 180
rect 485 145 500 165
rect 525 170 540 430
rect 565 240 580 465
rect 835 510 850 525
rect 835 475 885 485
rect 835 455 855 475
rect 875 455 885 475
rect 835 445 885 455
rect 835 425 850 445
rect 765 355 780 375
rect 835 365 850 375
rect 725 340 780 355
rect 805 350 850 365
rect 725 320 740 340
rect 725 245 740 270
rect 565 230 605 240
rect 565 210 575 230
rect 595 215 605 230
rect 700 235 740 245
rect 700 215 710 235
rect 730 215 740 235
rect 595 210 645 215
rect 565 200 645 210
rect 700 205 740 215
rect 525 155 570 170
rect 555 145 570 155
rect 555 75 570 95
rect 555 65 605 75
rect 555 45 575 65
rect 595 45 605 65
rect 555 35 605 45
rect 555 -5 570 10
rect 485 -70 500 -55
rect 555 -65 570 -55
rect 630 -65 645 200
rect 725 180 740 205
rect 725 115 740 130
rect 805 90 820 350
rect 910 320 925 585
rect 725 80 820 90
rect 725 60 735 80
rect 755 75 820 80
rect 845 310 925 320
rect 845 290 855 310
rect 875 305 925 310
rect 875 290 885 305
rect 845 280 885 290
rect 755 60 765 75
rect 725 50 765 60
rect 845 55 860 280
rect 725 30 740 50
rect 845 40 885 55
rect 870 30 885 40
rect 725 -35 740 -20
rect 870 -40 885 -20
rect 555 -80 645 -65
rect 845 -50 885 -40
rect 845 -70 855 -50
rect 875 -70 885 -50
rect 845 -80 885 -70
<< polycont >>
rect 575 570 595 590
rect 455 440 475 460
rect 430 285 450 305
rect 855 455 875 475
rect 575 210 595 230
rect 710 215 730 235
rect 575 45 595 65
rect 735 60 755 80
rect 855 290 875 310
rect 855 -70 875 -50
<< locali >>
rect 565 590 605 600
rect 565 580 575 590
rect 420 570 575 580
rect 595 570 605 590
rect 420 560 605 570
rect 680 565 760 575
rect 680 560 730 565
rect 420 540 440 560
rect 400 525 440 540
rect 400 505 410 525
rect 430 505 440 525
rect 400 490 440 505
rect 465 525 585 540
rect 465 505 475 525
rect 495 505 515 525
rect 535 505 555 525
rect 575 505 585 525
rect 465 490 585 505
rect 610 525 650 540
rect 610 505 620 525
rect 640 505 650 525
rect 610 490 650 505
rect 445 460 485 470
rect 445 440 455 460
rect 475 440 485 460
rect 445 430 485 440
rect 465 390 485 430
rect 400 375 440 390
rect 400 355 410 375
rect 430 355 440 375
rect 400 340 440 355
rect 465 375 505 390
rect 465 355 475 375
rect 495 360 505 375
rect 610 360 630 490
rect 680 390 690 560
rect 710 390 730 560
rect 680 380 730 390
rect 750 380 760 565
rect 680 375 760 380
rect 785 565 825 575
rect 785 380 795 565
rect 815 380 825 565
rect 855 560 895 575
rect 855 540 865 560
rect 885 540 895 560
rect 855 525 895 540
rect 865 485 885 525
rect 845 475 885 485
rect 845 455 855 475
rect 875 455 885 475
rect 845 445 885 455
rect 785 375 825 380
rect 855 410 895 425
rect 855 390 865 410
rect 885 390 895 410
rect 855 375 895 390
rect 495 355 670 360
rect 465 340 670 355
rect 650 320 670 340
rect 855 320 875 375
rect 420 305 460 315
rect 400 285 430 305
rect 450 295 460 305
rect 650 305 720 320
rect 650 300 690 305
rect 450 285 630 295
rect 420 280 630 285
rect 680 285 690 300
rect 710 285 720 305
rect 420 275 645 280
rect 610 260 645 275
rect 680 270 720 285
rect 745 310 930 320
rect 745 305 855 310
rect 745 285 755 305
rect 775 300 855 305
rect 775 285 785 300
rect 745 270 785 285
rect 845 290 855 300
rect 875 300 930 310
rect 875 290 885 300
rect 845 280 885 290
rect 400 235 440 250
rect 400 215 410 235
rect 430 215 440 235
rect 400 200 440 215
rect 465 235 505 250
rect 625 245 645 260
rect 465 215 475 235
rect 495 220 505 235
rect 565 230 605 240
rect 565 220 575 230
rect 495 215 575 220
rect 465 210 575 215
rect 595 210 605 230
rect 625 235 930 245
rect 625 225 710 235
rect 465 200 605 210
rect 700 215 710 225
rect 730 225 930 235
rect 730 215 740 225
rect 700 205 740 215
rect 575 180 670 200
rect 575 145 595 180
rect 650 165 720 180
rect 650 160 690 165
rect 680 145 690 160
rect 710 145 720 165
rect 400 135 480 145
rect 400 130 450 135
rect 400 -40 410 130
rect 430 -40 450 130
rect 400 -45 450 -40
rect 470 -45 480 135
rect 400 -55 480 -45
rect 505 135 545 145
rect 505 -45 515 135
rect 535 -45 545 135
rect 575 130 615 145
rect 680 130 720 145
rect 745 165 930 180
rect 745 145 755 165
rect 775 160 930 165
rect 775 145 785 160
rect 745 130 785 145
rect 575 110 585 130
rect 605 110 615 130
rect 575 95 615 110
rect 745 90 765 130
rect 725 80 765 90
rect 565 65 605 75
rect 565 45 575 65
rect 595 45 605 65
rect 725 60 735 80
rect 755 60 765 80
rect 725 50 765 60
rect 565 35 605 45
rect 585 -5 605 35
rect 890 30 910 160
rect 680 15 720 30
rect 680 -5 690 15
rect 710 -5 720 15
rect 505 -55 545 -45
rect 575 -20 615 -5
rect 680 -20 720 -5
rect 745 15 865 30
rect 745 -5 755 15
rect 775 -5 795 15
rect 815 -5 835 15
rect 855 -5 865 15
rect 745 -20 865 -5
rect 890 15 930 30
rect 890 -5 900 15
rect 920 -5 930 15
rect 890 -20 930 -5
rect 575 -40 585 -20
rect 605 -40 615 -20
rect 575 -55 615 -40
rect 700 -40 720 -20
rect 700 -50 885 -40
rect 700 -60 855 -50
rect 845 -70 855 -60
rect 875 -70 885 -50
rect 845 -80 885 -70
<< viali >>
rect 515 505 535 525
rect 690 390 710 560
rect 410 -40 430 130
rect 795 -5 815 15
<< metal1 >>
rect -75 95 175 210
rect -75 -55 175 60
<< end >>
