* SPICE3 file created from m2m_ladder.ext - technology: sky130A

X0 a_8000_7800# a_5600_9530# IOUT VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X1 a_20600_7800# D2 IDUMP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X2 a_22600_9530# D1 VP VP sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X3 a_27000_9530# D0 VP VP sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X4 a_25000_13400# VGATE a_20600_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X5 a_12200_7800# a_9800_9530# IOUT VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X6 a_3800_13400# VGATE IIN VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X7 a_20600_13400# VGATE a_16400_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X8 a_25000_13400# VGATE a_20600_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X9 a_25000_7800# a_22600_9530# IOUT VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X10 a_29400_7800# a_27000_9530# IOUT VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X11 a_1400_9530# D6 VN VN sky130_fd_pr__nfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X12 a_9800_9530# D4 VP VP sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X13 a_3800_13400# VGATE IIN VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X14 a_20600_13400# VGATE a_16400_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X15 a_25000_7800# VGATE a_20600_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X16 a_3800_7800# VGATE IIN VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X17 a_20600_7800# VGATE a_16400_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X18 a_3800_7800# D6 IDUMP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X19 a_5600_9530# D5 VN VN sky130_fd_pr__nfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X20 a_14000_9530# D3 VP VP sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X21 a_16400_13400# VGATE a_12200_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X22 a_16400_13400# VGATE a_12200_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X23 a_16400_7800# a_14000_9530# IOUT VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X24 a_8000_7800# D5 IDUMP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X25 a_22600_9530# D1 VN VN sky130_fd_pr__nfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X26 a_27000_9530# D0 VN VN sky130_fd_pr__nfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X27 a_18200_9530# D2 VP VP sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X28 a_16400_7800# VGATE a_12200_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X29 a_29400_13400# VGATE a_25000_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=12 as=16 ps=16 w=4 l=12
X30 a_12200_13400# VGATE a_8000_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X31 a_29400_13400# VGATE a_25000_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=12 as=16 ps=16 w=4 l=12
X32 a_20600_7800# a_18200_9530# IOUT VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X33 a_12200_7800# D4 IDUMP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X34 a_25000_7800# D1 IDUMP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X35 a_29400_7800# D0 IDUMP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X36 a_9800_9530# D4 VN VN sky130_fd_pr__nfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X37 a_12200_13400# VGATE a_8000_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X38 a_29400_7800# VGATE a_25000_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X39 a_12200_7800# VGATE a_8000_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X40 a_1400_9530# D6 VP VP sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X41 a_14000_9530# D3 VN VN sky130_fd_pr__nfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X42 a_3800_7800# a_1400_9530# IOUT VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X43 a_8000_13400# VGATE a_3800_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X44 IDUMP VGATE a_29400_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=12 w=4 l=12
X45 a_5600_9530# D5 VP VP sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X46 a_8000_13400# VGATE a_3800_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X47 a_16400_7800# D3 IDUMP VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
X48 a_18200_9530# D2 VN VN sky130_fd_pr__nfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X49 IDUMP VGATE a_29400_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=12 w=4 l=12
X50 a_8000_7800# VGATE a_3800_13400# VP sky130_fd_pr__pfet_01v8 ad=16 pd=16 as=16 ps=16 w=4 l=12
