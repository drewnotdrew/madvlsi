* SPICE3 file created from shift_register.ext - technology: sky130A

X0 csrl_edge_0/a_1410_1020# clk VP VP sky130_fd_pr__pfet_01v8 ad=0.33332 pd=1.765 as=0.9 ps=4.9 w=2 l=0.15
X1 csrl_edge_0/a_1000_n110# clk VN VN sky130_fd_pr__nfet_01v8 ad=0.33332 pd=1.765 as=0.9 ps=4.9 w=2 l=0.15
X2 VN csrl_edge_1/Dn csrl_edge_1/D VN sky130_fd_pr__nfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X3 csrl_edge_1/D clk csrl_edge_0/a_800_1290# VN sky130_fd_pr__nfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X4 csrl_edge_0/a_800_980# csrl_edge_0/a_800_1290# csrl_edge_0/a_1000_n110# VN sky130_fd_pr__nfet_01v8 ad=0.225 pd=1.9 as=0.33332 ps=1.765 w=0.5 l=0.15
X5 VP csrl_edge_0/a_800_980# csrl_edge_0/a_800_1290# VP sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X6 csrl_edge_0/a_800_1290# csrl_edge_0/a_800_980# csrl_edge_0/a_1000_n110# VN sky130_fd_pr__nfet_01v8 ad=0.225 pd=1.9 as=0.33332 ps=1.765 w=0.5 l=0.15
X7 csrl_edge_1/D csrl_edge_1/Dn csrl_edge_0/a_1410_1020# VP sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.9 as=0.33332 ps=1.765 w=0.5 l=0.15
X8 csrl_edge_1/Dn csrl_edge_1/D csrl_edge_0/a_1410_1020# VP sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.9 as=0.33332 ps=1.765 w=0.5 l=0.15
X9 csrl_edge_1/Dn clk csrl_edge_0/a_800_980# VN sky130_fd_pr__nfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X10 VN csrl_edge_1/D csrl_edge_1/Dn VN sky130_fd_pr__nfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X11 csrl_edge_0/a_800_1290# clk D VP sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X12 VP csrl_edge_0/a_800_1290# csrl_edge_0/a_800_980# VP sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X13 csrl_edge_0/a_800_980# clk Dn VP sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.9 as=0.225 ps=1.9 w=0.5 l=0.15
X14 csrl_edge_1/a_1410_1020# clk VP VP sky130_fd_pr__pfet_01v8 ad=1 pd=5.3 as=5.4 ps=34.8 w=2 l=0.15
X15 csrl_edge_1/a_1000_n110# clk VN VN sky130_fd_pr__nfet_01v8 ad=1 pd=5.3 as=5.4 ps=34.8 w=2 l=0.15
X16 VN csrl_edge_2/Dn csrl_edge_2/D VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.45 ps=3.8 w=0.5 l=0.15
X17 csrl_edge_2/D clk csrl_edge_1/a_800_1290# VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.45 ps=3.8 w=0.5 l=0.15
X18 csrl_edge_1/a_800_980# csrl_edge_1/a_800_1290# csrl_edge_1/a_1000_n110# VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=3.8 as=0 ps=0 w=0.5 l=0.15
X19 VP csrl_edge_1/a_800_980# csrl_edge_1/a_800_1290# VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.45 ps=3.8 w=0.5 l=0.15
X20 csrl_edge_1/a_800_1290# csrl_edge_1/a_800_980# csrl_edge_1/a_1000_n110# VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.15
X21 csrl_edge_2/D csrl_edge_2/Dn csrl_edge_1/a_1410_1020# VP sky130_fd_pr__pfet_01v8 ad=0.45 pd=3.8 as=0 ps=0 w=0.5 l=0.15
X22 csrl_edge_2/Dn csrl_edge_2/D csrl_edge_1/a_1410_1020# VP sky130_fd_pr__pfet_01v8 ad=0.45 pd=3.8 as=0 ps=0 w=0.5 l=0.15
X23 csrl_edge_2/Dn clk csrl_edge_1/a_800_980# VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=3.8 as=0 ps=0 w=0.5 l=0.15
X24 VN csrl_edge_2/D csrl_edge_2/Dn VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.15
X25 csrl_edge_1/a_800_1290# clk csrl_edge_1/D VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.45 ps=3.8 w=0.5 l=0.15
X26 VP csrl_edge_1/a_800_1290# csrl_edge_1/a_800_980# VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.45 ps=3.8 w=0.5 l=0.15
X27 csrl_edge_1/a_800_980# clk csrl_edge_1/Dn VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.45 ps=3.8 w=0.5 l=0.15
X28 csrl_edge_2/a_1410_1020# clk VP VP sky130_fd_pr__pfet_01v8 ad=1 pd=5.3 as=0 ps=0 w=2 l=0.15
X29 csrl_edge_2/a_1000_n110# clk VN VN sky130_fd_pr__nfet_01v8 ad=1 pd=5.3 as=0 ps=0 w=2 l=0.15
X30 VN csrl_edge_3/Dn csrl_edge_3/D VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.45 ps=3.8 w=0.5 l=0.15
X31 csrl_edge_3/D clk csrl_edge_2/a_800_1290# VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.45 ps=3.8 w=0.5 l=0.15
X32 csrl_edge_2/a_800_980# csrl_edge_2/a_800_1290# csrl_edge_2/a_1000_n110# VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=3.8 as=0 ps=0 w=0.5 l=0.15
X33 VP csrl_edge_2/a_800_980# csrl_edge_2/a_800_1290# VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.45 ps=3.8 w=0.5 l=0.15
X34 csrl_edge_2/a_800_1290# csrl_edge_2/a_800_980# csrl_edge_2/a_1000_n110# VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.15
X35 csrl_edge_3/D csrl_edge_3/Dn csrl_edge_2/a_1410_1020# VP sky130_fd_pr__pfet_01v8 ad=0.45 pd=3.8 as=0 ps=0 w=0.5 l=0.15
X36 csrl_edge_3/Dn csrl_edge_3/D csrl_edge_2/a_1410_1020# VP sky130_fd_pr__pfet_01v8 ad=0.45 pd=3.8 as=0 ps=0 w=0.5 l=0.15
X37 csrl_edge_3/Dn clk csrl_edge_2/a_800_980# VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=3.8 as=0 ps=0 w=0.5 l=0.15
X38 VN csrl_edge_3/D csrl_edge_3/Dn VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.15
X39 csrl_edge_2/a_800_1290# clk csrl_edge_2/D VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.15
X40 VP csrl_edge_2/a_800_1290# csrl_edge_2/a_800_980# VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.45 ps=3.8 w=0.5 l=0.15
X41 csrl_edge_2/a_800_980# clk csrl_edge_2/Dn VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.15
X42 csrl_edge_3/a_1410_1020# clk VP VP sky130_fd_pr__pfet_01v8 ad=1 pd=5.3 as=0 ps=0 w=2 l=0.15
X43 csrl_edge_3/a_1000_n110# clk VN VN sky130_fd_pr__nfet_01v8 ad=1 pd=5.3 as=0 ps=0 w=2 l=0.15
X44 VN Qn Q VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.45 ps=3.8 w=0.5 l=0.15
X45 Q clk csrl_edge_3/a_800_1290# VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.45 ps=3.8 w=0.5 l=0.15
X46 csrl_edge_3/a_800_980# csrl_edge_3/a_800_1290# csrl_edge_3/a_1000_n110# VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=3.8 as=0 ps=0 w=0.5 l=0.15
X47 VP csrl_edge_3/a_800_980# csrl_edge_3/a_800_1290# VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.45 ps=3.8 w=0.5 l=0.15
X48 csrl_edge_3/a_800_1290# csrl_edge_3/a_800_980# csrl_edge_3/a_1000_n110# VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.15
X49 Q Qn csrl_edge_3/a_1410_1020# VP sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.9 as=0 ps=0 w=0.5 l=0.15
X50 Qn Q csrl_edge_3/a_1410_1020# VP sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.9 as=0 ps=0 w=0.5 l=0.15
X51 Qn clk csrl_edge_3/a_800_980# VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=3.8 as=0 ps=0 w=0.5 l=0.15
X52 VN Q Qn VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.15
X53 csrl_edge_3/a_800_1290# clk csrl_edge_3/D VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.15
X54 VP csrl_edge_3/a_800_1290# csrl_edge_3/a_800_980# VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.45 ps=3.8 w=0.5 l=0.15
X55 csrl_edge_3/a_800_980# clk csrl_edge_3/Dn VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.15
