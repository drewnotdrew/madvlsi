** sch_path: /home/drew/Documents/git/madvlsi/dac/schematic/m2m_ladder_tb.sch
**.subckt m2m_ladder_tb
Vb0 b0 GND 1
Vb1 b1 GND 1
Vb2 b2 GND 1
Vb3 b3 GND 1
Vb4 b4 GND 1
Vb5 b5 GND 1
Vb6 b6 GND 1
I1 GND I_in 1m
V1 V_gate GND 1
V2 VDD GND 1.8
Vout net1 GND 0
.save i(vout)
**** begin user architecture code


.control
  set wr_vecnames
  set wr_singlescale
  let code = 0
  while code < 128
    if code eq 0
      let b0 = 0
    else
      let b0 = code % 2
    end
    if floor(code / 2) eq 0
      let b1 = 0
    else
      let b1 = floor(code / 2) % 2
    end
    if floor(code / 4) eq 0
      let b2 = 0
    else
      let b2 = floor(code / 4) % 2
    end
    if floor(code / 8) eq 0
      let b3 = 0
    else
      let b3 = floor(code / 8) % 2
    end
    if floor(code / 16) eq 0
      let b4 = 0
    else
      let b4 = floor(code / 16) % 2
    end
    if floor(code / 32) eq 0
      let b5 = 0
    else
      let b5 = floor(code / 32) % 2
    end
    if floor(code / 64) eq 0
      let b6 = 0
    else
      let b6 = floor(code / 64) % 2
    end
    alter vb0 $&b0
    alter vb1 $&b1
    alter vb2 $&b2
    alter vb3 $&b3
    alter vb4 $&b4
    alter vb5 $&b5
    alter vb6 $&b6
    save all
    op
    wrdata ~/documents/git/madvlsi/dac/schematic/m2m_ladder_tb.txt v(b0) v(b1) v(b2) v(b3) v(b4) v(b5) v(b6) i(Vout)
    if code eq 0
      set appendwrite
      set wr_vecnames = FALSE
    end
    let code = code + 1
  end
  quit
.endc

.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt
**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
