magic
tech sky130A
timestamp 1763181149
<< nwell >>
rect 250 6200 17150 8100
rect 250 3700 15600 6200
rect 250 2700 1200 3700
rect 1495 3500 3300 3700
rect 3595 3500 5400 3700
rect 5695 3500 7500 3700
rect 7795 3500 9600 3700
rect 9995 3500 11800 3700
rect 12195 3500 14000 3700
rect 14395 3500 15600 3700
rect 1500 2700 3300 3500
rect 3600 2700 5400 3500
rect 5700 2700 7500 3500
rect 7800 2700 9600 3500
rect 10000 2700 11800 3500
rect 12200 2700 14000 3500
rect 14400 2700 15600 3500
<< nmos >>
rect 1340 3575 1355 3625
rect 3440 3575 3455 3625
rect 5540 3575 5555 3625
rect 7640 3575 7655 3625
rect 9740 3575 9755 3625
rect 11940 3575 11955 3625
rect 14140 3575 14155 3625
<< pmos >>
rect 700 7200 1900 7600
rect 2800 7200 4000 7600
rect 4900 7200 6100 7600
rect 7000 7200 8200 7600
rect 9100 7200 10300 7600
rect 11300 7200 12500 7600
rect 13500 7200 14700 7600
rect 15500 7200 16700 7600
rect 700 6700 1900 7100
rect 2800 6700 4000 7100
rect 4900 6700 6100 7100
rect 7000 6700 8200 7100
rect 9100 6700 10300 7100
rect 11300 6700 12500 7100
rect 13500 6700 14700 7100
rect 15500 6700 16700 7100
rect 700 5700 1900 6100
rect 2800 5700 4000 6100
rect 4900 5700 6100 6100
rect 7000 5700 8200 6100
rect 9100 5700 10300 6100
rect 11300 5700 12500 6100
rect 13500 5700 14700 6100
rect 700 4800 1900 5200
rect 2800 4800 4000 5200
rect 4900 4800 6100 5200
rect 7000 4800 8200 5200
rect 9100 4800 10300 5200
rect 11300 4800 12500 5200
rect 13500 4800 14700 5200
rect 700 3900 1900 4300
rect 2800 3900 4000 4300
rect 4900 3900 6100 4300
rect 7000 3900 8200 4300
rect 9100 3900 10300 4300
rect 11300 3900 12500 4300
rect 13500 3900 14700 4300
rect 1340 3775 1355 3825
rect 3440 3775 3455 3825
rect 5540 3775 5555 3825
rect 7640 3775 7655 3825
rect 9740 3775 9755 3825
rect 11940 3775 11955 3825
rect 14140 3775 14155 3825
<< ndiff >>
rect 1295 3610 1340 3625
rect 1295 3590 1305 3610
rect 1325 3590 1340 3610
rect 1295 3575 1340 3590
rect 1355 3610 1400 3625
rect 1355 3590 1370 3610
rect 1390 3590 1400 3610
rect 1355 3575 1400 3590
rect 3395 3610 3440 3625
rect 3395 3590 3405 3610
rect 3425 3590 3440 3610
rect 3395 3575 3440 3590
rect 3455 3610 3500 3625
rect 3455 3590 3470 3610
rect 3490 3590 3500 3610
rect 3455 3575 3500 3590
rect 5495 3610 5540 3625
rect 5495 3590 5505 3610
rect 5525 3590 5540 3610
rect 5495 3575 5540 3590
rect 5555 3610 5600 3625
rect 5555 3590 5570 3610
rect 5590 3590 5600 3610
rect 5555 3575 5600 3590
rect 7595 3610 7640 3625
rect 7595 3590 7605 3610
rect 7625 3590 7640 3610
rect 7595 3575 7640 3590
rect 7655 3610 7700 3625
rect 7655 3590 7670 3610
rect 7690 3590 7700 3610
rect 7655 3575 7700 3590
rect 9695 3610 9740 3625
rect 9695 3590 9705 3610
rect 9725 3590 9740 3610
rect 9695 3575 9740 3590
rect 9755 3610 9800 3625
rect 9755 3590 9770 3610
rect 9790 3590 9800 3610
rect 9755 3575 9800 3590
rect 11895 3610 11940 3625
rect 11895 3590 11905 3610
rect 11925 3590 11940 3610
rect 11895 3575 11940 3590
rect 11955 3610 12000 3625
rect 11955 3590 11970 3610
rect 11990 3590 12000 3610
rect 11955 3575 12000 3590
rect 14095 3610 14140 3625
rect 14095 3590 14105 3610
rect 14125 3590 14140 3610
rect 14095 3575 14140 3590
rect 14155 3610 14200 3625
rect 14155 3590 14170 3610
rect 14190 3590 14200 3610
rect 14155 3575 14200 3590
<< pdiff >>
rect 300 7500 700 7600
rect 300 7300 400 7500
rect 600 7300 700 7500
rect 300 7200 700 7300
rect 1900 7500 2300 7600
rect 1900 7300 2000 7500
rect 2200 7300 2300 7500
rect 1900 7200 2300 7300
rect 2400 7500 2800 7600
rect 2400 7300 2500 7500
rect 2700 7300 2800 7500
rect 2400 7200 2800 7300
rect 4000 7500 4400 7600
rect 4000 7300 4100 7500
rect 4300 7300 4400 7500
rect 4000 7200 4400 7300
rect 4500 7500 4900 7600
rect 4500 7300 4600 7500
rect 4800 7300 4900 7500
rect 4500 7200 4900 7300
rect 6100 7500 6500 7600
rect 6100 7300 6200 7500
rect 6400 7300 6500 7500
rect 6100 7200 6500 7300
rect 6600 7500 7000 7600
rect 6600 7300 6700 7500
rect 6900 7300 7000 7500
rect 6600 7200 7000 7300
rect 8200 7500 8600 7600
rect 8200 7300 8300 7500
rect 8500 7300 8600 7500
rect 8200 7200 8600 7300
rect 8700 7500 9100 7600
rect 8700 7300 8800 7500
rect 9000 7300 9100 7500
rect 8700 7200 9100 7300
rect 10300 7500 10700 7600
rect 10300 7300 10400 7500
rect 10600 7300 10700 7500
rect 10300 7200 10700 7300
rect 10900 7500 11300 7600
rect 10900 7300 11000 7500
rect 11200 7300 11300 7500
rect 10900 7200 11300 7300
rect 12500 7500 12900 7600
rect 12500 7300 12600 7500
rect 12800 7300 12900 7500
rect 12500 7200 12900 7300
rect 13100 7500 13500 7600
rect 13100 7300 13200 7500
rect 13400 7300 13500 7500
rect 13100 7200 13500 7300
rect 14700 7500 15500 7600
rect 14700 7300 14800 7500
rect 15000 7300 15200 7500
rect 15400 7300 15500 7500
rect 14700 7200 15500 7300
rect 16700 7500 17100 7600
rect 16700 7300 16800 7500
rect 17000 7300 17100 7500
rect 16700 7200 17100 7300
rect 300 7000 700 7100
rect 300 6800 400 7000
rect 600 6800 700 7000
rect 300 6700 700 6800
rect 1900 7000 2300 7100
rect 1900 6800 2000 7000
rect 2200 6800 2300 7000
rect 1900 6700 2300 6800
rect 2400 7000 2800 7100
rect 2400 6800 2500 7000
rect 2700 6800 2800 7000
rect 2400 6700 2800 6800
rect 4000 7000 4400 7100
rect 4000 6800 4100 7000
rect 4300 6800 4400 7000
rect 4000 6700 4400 6800
rect 4500 7000 4900 7100
rect 4500 6800 4600 7000
rect 4800 6800 4900 7000
rect 4500 6700 4900 6800
rect 6100 7000 6500 7100
rect 6100 6800 6200 7000
rect 6400 6800 6500 7000
rect 6100 6700 6500 6800
rect 6600 7000 7000 7100
rect 6600 6800 6700 7000
rect 6900 6800 7000 7000
rect 6600 6700 7000 6800
rect 8200 7000 8600 7100
rect 8200 6800 8300 7000
rect 8500 6800 8600 7000
rect 8200 6700 8600 6800
rect 8700 7000 9100 7100
rect 8700 6800 8800 7000
rect 9000 6800 9100 7000
rect 8700 6700 9100 6800
rect 10300 7000 10700 7100
rect 10300 6800 10400 7000
rect 10600 6800 10700 7000
rect 10300 6700 10700 6800
rect 10900 7000 11300 7100
rect 10900 6800 11000 7000
rect 11200 6800 11300 7000
rect 10900 6700 11300 6800
rect 12500 7000 12900 7100
rect 12500 6800 12600 7000
rect 12800 6800 12900 7000
rect 12500 6700 12900 6800
rect 13100 7000 13500 7100
rect 13100 6800 13200 7000
rect 13400 6800 13500 7000
rect 13100 6700 13500 6800
rect 14700 7000 15500 7100
rect 14700 6800 14800 7000
rect 15000 6800 15200 7000
rect 15400 6800 15500 7000
rect 14700 6700 15500 6800
rect 16700 7000 17100 7100
rect 16700 6800 16800 7000
rect 17000 6800 17100 7000
rect 16700 6700 17100 6800
rect 300 6000 700 6100
rect 300 5800 400 6000
rect 600 5800 700 6000
rect 300 5700 700 5800
rect 1900 6000 2300 6100
rect 1900 5800 2000 6000
rect 2200 5800 2300 6000
rect 1900 5700 2300 5800
rect 2400 6000 2800 6100
rect 2400 5800 2500 6000
rect 2700 5800 2800 6000
rect 2400 5700 2800 5800
rect 4000 6000 4400 6100
rect 4000 5800 4100 6000
rect 4300 5800 4400 6000
rect 4000 5700 4400 5800
rect 4500 6000 4900 6100
rect 4500 5800 4600 6000
rect 4800 5800 4900 6000
rect 4500 5700 4900 5800
rect 6100 6000 6500 6100
rect 6100 5800 6200 6000
rect 6400 5800 6500 6000
rect 6100 5700 6500 5800
rect 6600 6000 7000 6100
rect 6600 5800 6700 6000
rect 6900 5800 7000 6000
rect 6600 5700 7000 5800
rect 8200 6000 8600 6100
rect 8200 5800 8300 6000
rect 8500 5800 8600 6000
rect 8200 5700 8600 5800
rect 8700 6000 9100 6100
rect 8700 5800 8800 6000
rect 9000 5800 9100 6000
rect 8700 5700 9100 5800
rect 10300 6000 10700 6100
rect 10300 5800 10400 6000
rect 10600 5800 10700 6000
rect 10300 5700 10700 5800
rect 10900 6000 11300 6100
rect 10900 5800 11000 6000
rect 11200 5800 11300 6000
rect 10900 5700 11300 5800
rect 12500 6000 12900 6100
rect 12500 5800 12600 6000
rect 12800 5800 12900 6000
rect 12500 5700 12900 5800
rect 13100 6000 13500 6100
rect 13100 5800 13200 6000
rect 13400 5800 13500 6000
rect 13100 5700 13500 5800
rect 14700 6000 15100 6100
rect 14700 5800 14800 6000
rect 15000 5800 15100 6000
rect 14700 5700 15100 5800
rect 300 5100 700 5200
rect 300 4900 400 5100
rect 600 4900 700 5100
rect 300 4800 700 4900
rect 1900 5100 2300 5200
rect 1900 4900 2000 5100
rect 2200 4900 2300 5100
rect 1900 4800 2300 4900
rect 2400 5100 2800 5200
rect 2400 4900 2500 5100
rect 2700 4900 2800 5100
rect 2400 4800 2800 4900
rect 4000 5100 4400 5200
rect 4000 4900 4100 5100
rect 4300 4900 4400 5100
rect 4000 4800 4400 4900
rect 4500 5100 4900 5200
rect 4500 4900 4600 5100
rect 4800 4900 4900 5100
rect 4500 4800 4900 4900
rect 6100 5100 6500 5200
rect 6100 4900 6200 5100
rect 6400 4900 6500 5100
rect 6100 4800 6500 4900
rect 6600 5100 7000 5200
rect 6600 4900 6700 5100
rect 6900 4900 7000 5100
rect 6600 4800 7000 4900
rect 8200 5100 8600 5200
rect 8200 4900 8300 5100
rect 8500 4900 8600 5100
rect 8200 4800 8600 4900
rect 8700 5100 9100 5200
rect 8700 4900 8800 5100
rect 9000 4900 9100 5100
rect 8700 4800 9100 4900
rect 10300 5100 10700 5200
rect 10300 4900 10400 5100
rect 10600 4900 10700 5100
rect 10300 4800 10700 4900
rect 10900 5100 11300 5200
rect 10900 4900 11000 5100
rect 11200 4900 11300 5100
rect 10900 4800 11300 4900
rect 12500 5100 12900 5200
rect 12500 4900 12600 5100
rect 12800 4900 12900 5100
rect 12500 4800 12900 4900
rect 13100 5100 13500 5200
rect 13100 4900 13200 5100
rect 13400 4900 13500 5100
rect 13100 4800 13500 4900
rect 14700 5100 15100 5200
rect 14700 4900 14800 5100
rect 15000 4900 15100 5100
rect 14700 4800 15100 4900
rect 300 4200 700 4300
rect 300 4000 400 4200
rect 600 4000 700 4200
rect 300 3900 700 4000
rect 1900 4200 2300 4300
rect 1900 4000 2000 4200
rect 2200 4000 2300 4200
rect 1900 3900 2300 4000
rect 2400 4200 2800 4300
rect 2400 4000 2500 4200
rect 2700 4000 2800 4200
rect 2400 3900 2800 4000
rect 4000 4200 4400 4300
rect 4000 4000 4100 4200
rect 4300 4000 4400 4200
rect 4000 3900 4400 4000
rect 4500 4200 4900 4300
rect 4500 4000 4600 4200
rect 4800 4000 4900 4200
rect 4500 3900 4900 4000
rect 6100 4200 6500 4300
rect 6100 4000 6200 4200
rect 6400 4000 6500 4200
rect 6100 3900 6500 4000
rect 6600 4200 7000 4300
rect 6600 4000 6700 4200
rect 6900 4000 7000 4200
rect 6600 3900 7000 4000
rect 8200 4200 8600 4300
rect 8200 4000 8300 4200
rect 8500 4000 8600 4200
rect 8200 3900 8600 4000
rect 8700 4200 9100 4300
rect 8700 4000 8800 4200
rect 9000 4000 9100 4200
rect 8700 3900 9100 4000
rect 10300 4200 10700 4300
rect 10300 4000 10400 4200
rect 10600 4000 10700 4200
rect 10300 3900 10700 4000
rect 10900 4200 11300 4300
rect 10900 4000 11000 4200
rect 11200 4000 11300 4200
rect 10900 3900 11300 4000
rect 12500 4200 12900 4300
rect 12500 4000 12600 4200
rect 12800 4000 12900 4200
rect 12500 3900 12900 4000
rect 13100 4200 13500 4300
rect 13100 4000 13200 4200
rect 13400 4000 13500 4200
rect 13100 3900 13500 4000
rect 14700 4200 15100 4300
rect 14700 4000 14800 4200
rect 15000 4000 15100 4200
rect 14700 3900 15100 4000
rect 1295 3810 1340 3825
rect 1295 3790 1305 3810
rect 1325 3790 1340 3810
rect 1295 3775 1340 3790
rect 1355 3810 1400 3825
rect 1355 3790 1370 3810
rect 1390 3790 1400 3810
rect 1355 3775 1400 3790
rect 3395 3810 3440 3825
rect 3395 3790 3405 3810
rect 3425 3790 3440 3810
rect 3395 3775 3440 3790
rect 3455 3810 3500 3825
rect 3455 3790 3470 3810
rect 3490 3790 3500 3810
rect 3455 3775 3500 3790
rect 5495 3810 5540 3825
rect 5495 3790 5505 3810
rect 5525 3790 5540 3810
rect 5495 3775 5540 3790
rect 5555 3810 5600 3825
rect 5555 3790 5570 3810
rect 5590 3790 5600 3810
rect 5555 3775 5600 3790
rect 7595 3810 7640 3825
rect 7595 3790 7605 3810
rect 7625 3790 7640 3810
rect 7595 3775 7640 3790
rect 7655 3810 7700 3825
rect 7655 3790 7670 3810
rect 7690 3790 7700 3810
rect 7655 3775 7700 3790
rect 9695 3810 9740 3825
rect 9695 3790 9705 3810
rect 9725 3790 9740 3810
rect 9695 3775 9740 3790
rect 9755 3810 9800 3825
rect 9755 3790 9770 3810
rect 9790 3790 9800 3810
rect 9755 3775 9800 3790
rect 11895 3810 11940 3825
rect 11895 3790 11905 3810
rect 11925 3790 11940 3810
rect 11895 3775 11940 3790
rect 11955 3810 12000 3825
rect 11955 3790 11970 3810
rect 11990 3790 12000 3810
rect 11955 3775 12000 3790
rect 14095 3810 14140 3825
rect 14095 3790 14105 3810
rect 14125 3790 14140 3810
rect 14095 3775 14140 3790
rect 14155 3810 14200 3825
rect 14155 3790 14170 3810
rect 14190 3790 14200 3810
rect 14155 3775 14200 3790
<< ndiffc >>
rect 1305 3590 1325 3610
rect 1370 3590 1390 3610
rect 3405 3590 3425 3610
rect 3470 3590 3490 3610
rect 5505 3590 5525 3610
rect 5570 3590 5590 3610
rect 7605 3590 7625 3610
rect 7670 3590 7690 3610
rect 9705 3590 9725 3610
rect 9770 3590 9790 3610
rect 11905 3590 11925 3610
rect 11970 3590 11990 3610
rect 14105 3590 14125 3610
rect 14170 3590 14190 3610
<< pdiffc >>
rect 400 7300 600 7500
rect 2000 7300 2200 7500
rect 2500 7300 2700 7500
rect 4100 7300 4300 7500
rect 4600 7300 4800 7500
rect 6200 7300 6400 7500
rect 6700 7300 6900 7500
rect 8300 7300 8500 7500
rect 8800 7300 9000 7500
rect 10400 7300 10600 7500
rect 11000 7300 11200 7500
rect 12600 7300 12800 7500
rect 13200 7300 13400 7500
rect 14800 7300 15000 7500
rect 15200 7300 15400 7500
rect 16800 7300 17000 7500
rect 400 6800 600 7000
rect 2000 6800 2200 7000
rect 2500 6800 2700 7000
rect 4100 6800 4300 7000
rect 4600 6800 4800 7000
rect 6200 6800 6400 7000
rect 6700 6800 6900 7000
rect 8300 6800 8500 7000
rect 8800 6800 9000 7000
rect 10400 6800 10600 7000
rect 11000 6800 11200 7000
rect 12600 6800 12800 7000
rect 13200 6800 13400 7000
rect 14800 6800 15000 7000
rect 15200 6800 15400 7000
rect 16800 6800 17000 7000
rect 400 5800 600 6000
rect 2000 5800 2200 6000
rect 2500 5800 2700 6000
rect 4100 5800 4300 6000
rect 4600 5800 4800 6000
rect 6200 5800 6400 6000
rect 6700 5800 6900 6000
rect 8300 5800 8500 6000
rect 8800 5800 9000 6000
rect 10400 5800 10600 6000
rect 11000 5800 11200 6000
rect 12600 5800 12800 6000
rect 13200 5800 13400 6000
rect 14800 5800 15000 6000
rect 400 4900 600 5100
rect 2000 4900 2200 5100
rect 2500 4900 2700 5100
rect 4100 4900 4300 5100
rect 4600 4900 4800 5100
rect 6200 4900 6400 5100
rect 6700 4900 6900 5100
rect 8300 4900 8500 5100
rect 8800 4900 9000 5100
rect 10400 4900 10600 5100
rect 11000 4900 11200 5100
rect 12600 4900 12800 5100
rect 13200 4900 13400 5100
rect 14800 4900 15000 5100
rect 400 4000 600 4200
rect 2000 4000 2200 4200
rect 2500 4000 2700 4200
rect 4100 4000 4300 4200
rect 4600 4000 4800 4200
rect 6200 4000 6400 4200
rect 6700 4000 6900 4200
rect 8300 4000 8500 4200
rect 8800 4000 9000 4200
rect 10400 4000 10600 4200
rect 11000 4000 11200 4200
rect 12600 4000 12800 4200
rect 13200 4000 13400 4200
rect 14800 4000 15000 4200
rect 1305 3790 1325 3810
rect 1370 3790 1390 3810
rect 3405 3790 3425 3810
rect 3470 3790 3490 3810
rect 5505 3790 5525 3810
rect 5570 3790 5590 3810
rect 7605 3790 7625 3810
rect 7670 3790 7690 3810
rect 9705 3790 9725 3810
rect 9770 3790 9790 3810
rect 11905 3790 11925 3810
rect 11970 3790 11990 3810
rect 14105 3790 14125 3810
rect 14170 3790 14190 3810
<< psubdiff >>
rect 1295 3435 1335 3450
rect 1295 3415 1305 3435
rect 1325 3415 1335 3435
rect 1295 3400 1335 3415
rect 3395 3435 3435 3450
rect 3395 3415 3405 3435
rect 3425 3415 3435 3435
rect 3395 3400 3435 3415
rect 5495 3435 5535 3450
rect 5495 3415 5505 3435
rect 5525 3415 5535 3435
rect 5495 3400 5535 3415
rect 7595 3435 7635 3450
rect 7595 3415 7605 3435
rect 7625 3415 7635 3435
rect 7595 3400 7635 3415
rect 9695 3435 9735 3450
rect 9695 3415 9705 3435
rect 9725 3415 9735 3435
rect 9695 3400 9735 3415
rect 11895 3435 11935 3450
rect 11895 3415 11905 3435
rect 11925 3415 11935 3435
rect 11895 3400 11935 3415
rect 14095 3435 14135 3450
rect 14095 3415 14105 3435
rect 14125 3415 14135 3435
rect 14095 3400 14135 3415
<< nsubdiff >>
rect 300 7950 700 8050
rect 300 7750 400 7950
rect 600 7750 700 7950
rect 300 7650 700 7750
rect 2200 7950 2600 8050
rect 2200 7750 2300 7950
rect 2500 7750 2600 7950
rect 2200 7650 2600 7750
rect 4300 7950 4700 8050
rect 4300 7750 4400 7950
rect 4600 7750 4700 7950
rect 4300 7650 4700 7750
rect 6400 7950 6800 8050
rect 6400 7750 6500 7950
rect 6700 7750 6800 7950
rect 6400 7650 6800 7750
rect 8500 7950 8900 8050
rect 8500 7750 8600 7950
rect 8800 7750 8900 7950
rect 8500 7650 8900 7750
rect 10600 7950 11000 8050
rect 10600 7750 10700 7950
rect 10900 7750 11000 7950
rect 10600 7650 11000 7750
rect 12800 7950 13200 8050
rect 12800 7750 12900 7950
rect 13100 7750 13200 7950
rect 12800 7650 13200 7750
rect 14900 7950 15300 8050
rect 14900 7750 15000 7950
rect 15200 7750 15300 7950
rect 14900 7650 15300 7750
rect 16700 7950 17100 8050
rect 16700 7750 16800 7950
rect 17000 7750 17100 7950
rect 16700 7650 17100 7750
rect 300 5550 700 5650
rect 300 5350 400 5550
rect 600 5350 700 5550
rect 300 5250 700 5350
rect 2400 5550 2800 5650
rect 2400 5350 2500 5550
rect 2700 5350 2800 5550
rect 2400 5250 2800 5350
rect 4500 5550 4900 5650
rect 4500 5350 4600 5550
rect 4800 5350 4900 5550
rect 4500 5250 4900 5350
rect 6600 5550 7000 5650
rect 6600 5350 6700 5550
rect 6900 5350 7000 5550
rect 6600 5250 7000 5350
rect 8700 5550 9100 5650
rect 8700 5350 8800 5550
rect 9000 5350 9100 5550
rect 8700 5250 9100 5350
rect 10900 5550 11300 5650
rect 10900 5350 11000 5550
rect 11200 5350 11300 5550
rect 10900 5250 11300 5350
rect 13100 5550 13500 5650
rect 13100 5350 13200 5550
rect 13400 5350 13500 5550
rect 13100 5250 13500 5350
rect 15150 5550 15550 5650
rect 15150 5350 15250 5550
rect 15450 5350 15550 5550
rect 15150 5250 15550 5350
rect 1225 3810 1265 3825
rect 1225 3790 1235 3810
rect 1255 3790 1265 3810
rect 1225 3775 1265 3790
rect 3325 3810 3365 3825
rect 3325 3790 3335 3810
rect 3355 3790 3365 3810
rect 3325 3775 3365 3790
rect 5425 3810 5465 3825
rect 5425 3790 5435 3810
rect 5455 3790 5465 3810
rect 5425 3775 5465 3790
rect 7525 3810 7565 3825
rect 7525 3790 7535 3810
rect 7555 3790 7565 3810
rect 7525 3775 7565 3790
rect 9625 3810 9665 3825
rect 9625 3790 9635 3810
rect 9655 3790 9665 3810
rect 9625 3775 9665 3790
rect 11825 3810 11865 3825
rect 11825 3790 11835 3810
rect 11855 3790 11865 3810
rect 11825 3775 11865 3790
rect 14025 3810 14065 3825
rect 14025 3790 14035 3810
rect 14055 3790 14065 3810
rect 14025 3775 14065 3790
rect 300 3200 700 3300
rect 300 3000 400 3200
rect 600 3000 700 3200
rect 300 2900 700 3000
rect 2400 3200 2800 3300
rect 2400 3000 2500 3200
rect 2700 3000 2800 3200
rect 2400 2900 2800 3000
rect 4500 3200 4900 3300
rect 4500 3000 4600 3200
rect 4800 3000 4900 3200
rect 4500 2900 4900 3000
rect 6600 3200 7000 3300
rect 6600 3000 6700 3200
rect 6900 3000 7000 3200
rect 6600 2900 7000 3000
rect 8700 3200 9100 3300
rect 8700 3000 8800 3200
rect 9000 3000 9100 3200
rect 8700 2900 9100 3000
rect 10900 3200 11300 3300
rect 10900 3000 11000 3200
rect 11200 3000 11300 3200
rect 10900 2900 11300 3000
rect 13100 3200 13500 3300
rect 13100 3000 13200 3200
rect 13400 3000 13500 3200
rect 13100 2900 13500 3000
rect 15150 3200 15550 3300
rect 15150 3000 15250 3200
rect 15450 3000 15550 3200
rect 15150 2900 15550 3000
<< psubdiffcont >>
rect 1305 3415 1325 3435
rect 3405 3415 3425 3435
rect 5505 3415 5525 3435
rect 7605 3415 7625 3435
rect 9705 3415 9725 3435
rect 11905 3415 11925 3435
rect 14105 3415 14125 3435
<< nsubdiffcont >>
rect 400 7750 600 7950
rect 2300 7750 2500 7950
rect 4400 7750 4600 7950
rect 6500 7750 6700 7950
rect 8600 7750 8800 7950
rect 10700 7750 10900 7950
rect 12900 7750 13100 7950
rect 15000 7750 15200 7950
rect 16800 7750 17000 7950
rect 400 5350 600 5550
rect 2500 5350 2700 5550
rect 4600 5350 4800 5550
rect 6700 5350 6900 5550
rect 8800 5350 9000 5550
rect 11000 5350 11200 5550
rect 13200 5350 13400 5550
rect 15250 5350 15450 5550
rect 1235 3790 1255 3810
rect 3335 3790 3355 3810
rect 5435 3790 5455 3810
rect 7535 3790 7555 3810
rect 9635 3790 9655 3810
rect 11835 3790 11855 3810
rect 14035 3790 14055 3810
rect 400 3000 600 3200
rect 2500 3000 2700 3200
rect 4600 3000 4800 3200
rect 6700 3000 6900 3200
rect 8800 3000 9000 3200
rect 11000 3000 11200 3200
rect 13200 3000 13400 3200
rect 15250 3000 15450 3200
<< poly >>
rect 700 7600 1900 7635
rect 2800 7600 4000 7635
rect 4900 7600 6100 7635
rect 7000 7600 8200 7635
rect 9100 7600 10300 7635
rect 11300 7600 12500 7635
rect 13500 7600 14700 7635
rect 15500 7600 16700 7635
rect 700 7100 1900 7200
rect 2800 7100 4000 7200
rect 4900 7100 6100 7200
rect 7000 7100 8200 7200
rect 9100 7100 10300 7200
rect 11300 7100 12500 7200
rect 13500 7100 14700 7200
rect 15500 7100 16700 7200
rect 700 6600 1900 6700
rect 2800 6600 4000 6700
rect 4900 6600 6100 6700
rect 7000 6600 8200 6700
rect 9100 6600 10300 6700
rect 11300 6600 12500 6700
rect 13500 6600 14700 6700
rect 15500 6600 16700 6700
rect -100 6200 16700 6600
rect 700 6100 1900 6200
rect 2800 6100 4000 6200
rect 4900 6100 6100 6200
rect 7000 6100 8200 6200
rect 9100 6100 10300 6200
rect 11300 6100 12500 6200
rect 13500 6100 14700 6200
rect 700 5665 1900 5700
rect 2800 5665 4000 5700
rect 4900 5665 6100 5700
rect 7000 5665 8200 5700
rect 9100 5665 10300 5700
rect 11300 5665 12500 5700
rect 13500 5665 14700 5700
rect 1400 5500 1800 5600
rect 1400 5300 1500 5500
rect 1700 5300 1800 5500
rect 1400 5235 1800 5300
rect 3500 5500 3900 5600
rect 3500 5300 3600 5500
rect 3800 5300 3900 5500
rect 3500 5235 3900 5300
rect 5600 5500 6000 5600
rect 5600 5300 5700 5500
rect 5900 5300 6000 5500
rect 5600 5235 6000 5300
rect 7700 5500 8100 5600
rect 7700 5300 7800 5500
rect 8000 5300 8100 5500
rect 7700 5235 8100 5300
rect 9800 5500 10200 5600
rect 9800 5300 9900 5500
rect 10100 5300 10200 5500
rect 9800 5235 10200 5300
rect 12000 5500 12400 5600
rect 12000 5300 12100 5500
rect 12300 5300 12400 5500
rect 12000 5235 12400 5300
rect 14200 5500 14600 5600
rect 14200 5300 14300 5500
rect 14500 5300 14600 5500
rect 14200 5235 14600 5300
rect 700 5200 1900 5235
rect 2800 5200 4000 5235
rect 4900 5200 6100 5235
rect 7000 5200 8200 5235
rect 9100 5200 10300 5235
rect 11300 5200 12500 5235
rect 13500 5200 14700 5235
rect 700 4765 1900 4800
rect 2800 4765 4000 4800
rect 4900 4765 6100 4800
rect 7000 4765 8200 4800
rect 9100 4765 10300 4800
rect 11300 4765 12500 4800
rect 13500 4765 14700 4800
rect 800 4600 1200 4700
rect 800 4400 900 4600
rect 1100 4400 1200 4600
rect 800 4335 1200 4400
rect 2900 4600 3300 4700
rect 2900 4400 3000 4600
rect 3200 4400 3300 4600
rect 2900 4335 3300 4400
rect 5000 4600 5400 4700
rect 5000 4400 5100 4600
rect 5300 4400 5400 4600
rect 5000 4335 5400 4400
rect 7100 4600 7500 4700
rect 7100 4400 7200 4600
rect 7400 4400 7500 4600
rect 7100 4335 7500 4400
rect 9200 4600 9600 4700
rect 9200 4400 9300 4600
rect 9500 4400 9600 4600
rect 9200 4335 9600 4400
rect 11400 4600 11800 4700
rect 11400 4400 11500 4600
rect 11700 4400 11800 4600
rect 11400 4335 11800 4400
rect 13600 4600 14000 4700
rect 13600 4400 13700 4600
rect 13900 4400 14000 4600
rect 13600 4335 14000 4400
rect 700 4300 1900 4335
rect 2800 4300 4000 4335
rect 4900 4300 6100 4335
rect 7000 4300 8200 4335
rect 9100 4300 10300 4335
rect 11300 4300 12500 4335
rect 13500 4300 14700 4335
rect 700 3865 1900 3900
rect 2800 3865 4000 3900
rect 4900 3865 6100 3900
rect 7000 3865 8200 3900
rect 9100 3865 10300 3900
rect 11300 3865 12500 3900
rect 13500 3865 14700 3900
rect 860 3800 1140 3840
rect 1340 3825 1355 3840
rect 860 3600 900 3800
rect 1100 3760 1140 3800
rect 2960 3800 3240 3840
rect 3440 3825 3455 3840
rect 1340 3760 1355 3775
rect 1100 3640 1355 3760
rect 1100 3600 1140 3640
rect 1340 3625 1355 3640
rect 860 3560 1140 3600
rect 2960 3600 3000 3800
rect 3200 3760 3240 3800
rect 5060 3800 5340 3840
rect 5540 3825 5555 3840
rect 3440 3760 3455 3775
rect 3200 3640 3455 3760
rect 3200 3600 3240 3640
rect 3440 3625 3455 3640
rect 1340 3560 1355 3575
rect 2960 3560 3240 3600
rect 5060 3600 5100 3800
rect 5300 3760 5340 3800
rect 7160 3800 7440 3840
rect 7640 3825 7655 3840
rect 5540 3760 5555 3775
rect 5300 3640 5555 3760
rect 5300 3600 5340 3640
rect 5540 3625 5555 3640
rect 3440 3560 3455 3575
rect 5060 3560 5340 3600
rect 7160 3600 7200 3800
rect 7400 3760 7440 3800
rect 9260 3800 9540 3840
rect 9740 3825 9755 3840
rect 7640 3760 7655 3775
rect 7400 3640 7655 3760
rect 7400 3600 7440 3640
rect 7640 3625 7655 3640
rect 5540 3560 5555 3575
rect 7160 3560 7440 3600
rect 9260 3600 9300 3800
rect 9500 3760 9540 3800
rect 11460 3800 11740 3840
rect 11940 3825 11955 3840
rect 9740 3760 9755 3775
rect 9500 3640 9755 3760
rect 9500 3600 9540 3640
rect 9740 3625 9755 3640
rect 7640 3560 7655 3575
rect 9260 3560 9540 3600
rect 11460 3600 11500 3800
rect 11700 3760 11740 3800
rect 13660 3800 13940 3840
rect 14140 3825 14155 3840
rect 11940 3760 11955 3775
rect 11700 3640 11955 3760
rect 11700 3600 11740 3640
rect 11940 3625 11955 3640
rect 9740 3560 9755 3575
rect 11460 3560 11740 3600
rect 13660 3600 13700 3800
rect 13900 3760 13940 3800
rect 14140 3760 14155 3775
rect 13900 3640 14155 3760
rect 13900 3600 13940 3640
rect 14140 3625 14155 3640
rect 11940 3560 11955 3575
rect 13660 3560 13940 3600
rect 14140 3560 14155 3575
<< polycont >>
rect 1500 5300 1700 5500
rect 3600 5300 3800 5500
rect 5700 5300 5900 5500
rect 7800 5300 8000 5500
rect 9900 5300 10100 5500
rect 12100 5300 12300 5500
rect 14300 5300 14500 5500
rect 900 4400 1100 4600
rect 3000 4400 3200 4600
rect 5100 4400 5300 4600
rect 7200 4400 7400 4600
rect 9300 4400 9500 4600
rect 11500 4400 11700 4600
rect 13700 4400 13900 4600
rect 900 3600 1100 3800
rect 3000 3600 3200 3800
rect 5100 3600 5300 3800
rect 7200 3600 7400 3800
rect 9300 3600 9500 3800
rect 11500 3600 11700 3800
rect 13700 3600 13900 3800
<< locali >>
rect 300 7950 700 8050
rect 300 7750 400 7950
rect 600 7750 700 7950
rect 300 7650 700 7750
rect 2200 7950 2600 8050
rect 2200 7750 2300 7950
rect 2500 7750 2600 7950
rect 2200 7650 2600 7750
rect 4300 7950 4700 8050
rect 4300 7750 4400 7950
rect 4600 7750 4700 7950
rect 4300 7650 4700 7750
rect 6400 7950 6800 8050
rect 6400 7750 6500 7950
rect 6700 7750 6800 7950
rect 6400 7650 6800 7750
rect 8500 7950 8900 8050
rect 8500 7750 8600 7950
rect 8800 7750 8900 7950
rect 8500 7650 8900 7750
rect 10600 7950 11000 8050
rect 10600 7750 10700 7950
rect 10900 7750 11000 7950
rect 10600 7650 11000 7750
rect 12800 7950 13200 8050
rect 12800 7750 12900 7950
rect 13100 7750 13200 7950
rect 12800 7650 13200 7750
rect 14900 7950 15300 8050
rect 14900 7750 15000 7950
rect 15200 7750 15300 7950
rect 14900 7650 15300 7750
rect 16700 7950 17100 8050
rect 16700 7750 16800 7950
rect 17000 7750 17100 7950
rect 16700 7650 17100 7750
rect 300 7500 700 7600
rect 300 7300 400 7500
rect 600 7300 700 7500
rect 300 7000 700 7300
rect 300 6800 400 7000
rect 600 6800 700 7000
rect 300 6600 700 6800
rect -50 6200 700 6600
rect 1900 7500 2300 7600
rect 1900 7300 2000 7500
rect 2200 7300 2300 7500
rect 1900 7000 2300 7300
rect 1900 6800 2000 7000
rect 2200 6800 2300 7000
rect 1900 6600 2300 6800
rect 2400 7500 2800 7600
rect 2400 7300 2500 7500
rect 2700 7300 2800 7500
rect 2400 7000 2800 7300
rect 2400 6800 2500 7000
rect 2700 6800 2800 7000
rect 2400 6600 2800 6800
rect 1900 6200 2800 6600
rect 4000 7500 4400 7600
rect 4000 7300 4100 7500
rect 4300 7300 4400 7500
rect 4000 7000 4400 7300
rect 4000 6800 4100 7000
rect 4300 6800 4400 7000
rect 4000 6600 4400 6800
rect 4500 7500 4900 7600
rect 4500 7300 4600 7500
rect 4800 7300 4900 7500
rect 4500 7000 4900 7300
rect 4500 6800 4600 7000
rect 4800 6800 4900 7000
rect 4500 6600 4900 6800
rect 4000 6200 4900 6600
rect 6100 7500 6500 7600
rect 6100 7300 6200 7500
rect 6400 7300 6500 7500
rect 6100 7000 6500 7300
rect 6100 6800 6200 7000
rect 6400 6800 6500 7000
rect 6100 6600 6500 6800
rect 6600 7500 7000 7600
rect 6600 7300 6700 7500
rect 6900 7300 7000 7500
rect 6600 7000 7000 7300
rect 6600 6800 6700 7000
rect 6900 6800 7000 7000
rect 6600 6600 7000 6800
rect 6100 6200 7000 6600
rect 8200 7500 8600 7600
rect 8200 7300 8300 7500
rect 8500 7300 8600 7500
rect 8200 7000 8600 7300
rect 8200 6800 8300 7000
rect 8500 6800 8600 7000
rect 8200 6600 8600 6800
rect 8700 7500 9100 7600
rect 8700 7300 8800 7500
rect 9000 7300 9100 7500
rect 8700 7000 9100 7300
rect 8700 6800 8800 7000
rect 9000 6800 9100 7000
rect 8700 6600 9100 6800
rect 8200 6200 9100 6600
rect 10300 7500 10700 7600
rect 10300 7300 10400 7500
rect 10600 7300 10700 7500
rect 10300 7000 10700 7300
rect 10300 6800 10400 7000
rect 10600 6800 10700 7000
rect 10300 6600 10700 6800
rect 10900 7500 11300 7600
rect 10900 7300 11000 7500
rect 11200 7300 11300 7500
rect 10900 7000 11300 7300
rect 10900 6800 11000 7000
rect 11200 6800 11300 7000
rect 10900 6600 11300 6800
rect 10300 6200 11300 6600
rect 12500 7500 12900 7600
rect 12500 7300 12600 7500
rect 12800 7300 12900 7500
rect 12500 7000 12900 7300
rect 12500 6800 12600 7000
rect 12800 6800 12900 7000
rect 12500 6600 12900 6800
rect 13100 7500 13500 7600
rect 13100 7300 13200 7500
rect 13400 7300 13500 7500
rect 13100 7000 13500 7300
rect 13100 6800 13200 7000
rect 13400 6800 13500 7000
rect 13100 6600 13500 6800
rect 14700 7500 15500 7600
rect 14700 7300 14800 7500
rect 15000 7300 15200 7500
rect 15400 7300 15500 7500
rect 14700 7000 15500 7300
rect 14700 6800 14800 7000
rect 15000 6800 15200 7000
rect 15400 6800 15500 7000
rect 14700 6700 15500 6800
rect 16700 7500 17100 7600
rect 16700 7300 16800 7500
rect 17000 7300 17100 7500
rect 16700 7000 17100 7300
rect 16700 6800 16800 7000
rect 17000 6800 17100 7000
rect 16700 6600 17100 6800
rect 12500 6200 13500 6600
rect 300 6000 700 6200
rect 300 5800 400 6000
rect 600 5800 700 6000
rect 300 5700 700 5800
rect 1900 6000 2300 6100
rect 1900 5800 2000 6000
rect 2200 5800 2300 6000
rect 300 5550 700 5650
rect 300 5350 400 5550
rect 600 5350 700 5550
rect 300 5250 700 5350
rect 1400 5500 1800 5600
rect 1400 5300 1500 5500
rect 1700 5300 1800 5500
rect 300 5100 700 5200
rect 300 4900 400 5100
rect 600 4900 700 5100
rect 300 4650 700 4900
rect 300 4450 400 4650
rect 600 4450 700 4650
rect 300 4350 700 4450
rect 800 4600 1200 4700
rect 800 4400 900 4600
rect 1100 4400 1200 4600
rect 300 4200 700 4300
rect 300 4000 400 4200
rect 600 4000 700 4200
rect 300 3800 700 4000
rect 300 3600 400 3800
rect 600 3600 700 3800
rect 300 3500 700 3600
rect 800 3800 1200 4400
rect 1400 3825 1800 5300
rect 1900 5100 2300 5800
rect 2400 6000 2800 6200
rect 2400 5800 2500 6000
rect 2700 5800 2800 6000
rect 2400 5700 2800 5800
rect 4000 6000 4400 6100
rect 4000 5800 4100 6000
rect 4300 5800 4400 6000
rect 2400 5550 2800 5650
rect 2400 5350 2500 5550
rect 2700 5350 2800 5550
rect 2400 5250 2800 5350
rect 3500 5500 3900 5600
rect 3500 5300 3600 5500
rect 3800 5300 3900 5500
rect 1900 4900 2000 5100
rect 2200 4900 2300 5100
rect 1900 4200 2300 4900
rect 2400 5100 2800 5200
rect 2400 4900 2500 5100
rect 2700 4900 2800 5100
rect 2400 4650 2800 4900
rect 2400 4450 2500 4650
rect 2700 4450 2800 4650
rect 2400 4350 2800 4450
rect 2900 4600 3300 4700
rect 2900 4400 3000 4600
rect 3200 4400 3300 4600
rect 1900 4000 2000 4200
rect 2200 4000 2300 4200
rect 1900 3900 2300 4000
rect 2400 4200 2800 4300
rect 2400 4000 2500 4200
rect 2700 4000 2800 4200
rect 800 3600 900 3800
rect 1100 3600 1200 3800
rect 800 3500 1200 3600
rect 1225 3810 1335 3825
rect 1225 3790 1235 3810
rect 1255 3790 1305 3810
rect 1325 3790 1335 3810
rect 1225 3775 1335 3790
rect 1360 3810 1800 3825
rect 1360 3790 1370 3810
rect 1390 3790 1800 3810
rect 300 3200 700 3300
rect 300 3000 400 3200
rect 600 3000 700 3200
rect 300 2900 700 3000
rect 900 2850 1100 3500
rect 1225 3290 1265 3775
rect 1295 3610 1335 3625
rect 1295 3590 1305 3610
rect 1325 3590 1335 3610
rect 1295 3435 1335 3590
rect 1360 3610 1800 3790
rect 1360 3590 1370 3610
rect 1390 3590 1800 3610
rect 1360 3575 1800 3590
rect 2400 3800 2800 4000
rect 2400 3600 2500 3800
rect 2700 3600 2800 3800
rect 2400 3500 2800 3600
rect 2900 3800 3300 4400
rect 3500 3825 3900 5300
rect 4000 5100 4400 5800
rect 4500 6000 4900 6200
rect 4500 5800 4600 6000
rect 4800 5800 4900 6000
rect 4500 5700 4900 5800
rect 6100 6000 6500 6100
rect 6100 5800 6200 6000
rect 6400 5800 6500 6000
rect 4500 5550 4900 5650
rect 4500 5350 4600 5550
rect 4800 5350 4900 5550
rect 4500 5250 4900 5350
rect 5600 5500 6000 5600
rect 5600 5300 5700 5500
rect 5900 5300 6000 5500
rect 4000 4900 4100 5100
rect 4300 4900 4400 5100
rect 4000 4200 4400 4900
rect 4500 5100 4900 5200
rect 4500 4900 4600 5100
rect 4800 4900 4900 5100
rect 4500 4650 4900 4900
rect 4500 4450 4600 4650
rect 4800 4450 4900 4650
rect 4500 4350 4900 4450
rect 5000 4600 5400 4700
rect 5000 4400 5100 4600
rect 5300 4400 5400 4600
rect 4000 4000 4100 4200
rect 4300 4000 4400 4200
rect 4000 3900 4400 4000
rect 4500 4200 4900 4300
rect 4500 4000 4600 4200
rect 4800 4000 4900 4200
rect 2900 3600 3000 3800
rect 3200 3600 3300 3800
rect 2900 3500 3300 3600
rect 3325 3810 3435 3825
rect 3325 3790 3335 3810
rect 3355 3790 3405 3810
rect 3425 3790 3435 3810
rect 3325 3775 3435 3790
rect 3460 3810 3900 3825
rect 3460 3790 3470 3810
rect 3490 3790 3900 3810
rect 1295 3415 1305 3435
rect 1325 3415 1335 3435
rect 1295 3400 1335 3415
rect 1225 3270 1235 3290
rect 1255 3270 1265 3290
rect 1225 3260 1265 3270
rect 2400 3200 2800 3300
rect 2400 3000 2500 3200
rect 2700 3000 2800 3200
rect 2400 2900 2800 3000
rect 3000 2850 3200 3500
rect 3325 3290 3365 3775
rect 3395 3610 3435 3625
rect 3395 3590 3405 3610
rect 3425 3590 3435 3610
rect 3395 3435 3435 3590
rect 3460 3610 3900 3790
rect 3460 3590 3470 3610
rect 3490 3590 3900 3610
rect 3460 3575 3900 3590
rect 4500 3800 4900 4000
rect 4500 3600 4600 3800
rect 4800 3600 4900 3800
rect 4500 3500 4900 3600
rect 5000 3800 5400 4400
rect 5600 3825 6000 5300
rect 6100 5100 6500 5800
rect 6600 6000 7000 6200
rect 6600 5800 6700 6000
rect 6900 5800 7000 6000
rect 6600 5700 7000 5800
rect 8200 6000 8600 6100
rect 8200 5800 8300 6000
rect 8500 5800 8600 6000
rect 6600 5550 7000 5650
rect 6600 5350 6700 5550
rect 6900 5350 7000 5550
rect 6600 5250 7000 5350
rect 7700 5500 8100 5600
rect 7700 5300 7800 5500
rect 8000 5300 8100 5500
rect 6100 4900 6200 5100
rect 6400 4900 6500 5100
rect 6100 4200 6500 4900
rect 6600 5100 7000 5200
rect 6600 4900 6700 5100
rect 6900 4900 7000 5100
rect 6600 4650 7000 4900
rect 6600 4450 6700 4650
rect 6900 4450 7000 4650
rect 6600 4350 7000 4450
rect 7100 4600 7500 4700
rect 7100 4400 7200 4600
rect 7400 4400 7500 4600
rect 6100 4000 6200 4200
rect 6400 4000 6500 4200
rect 6100 3900 6500 4000
rect 6600 4200 7000 4300
rect 6600 4000 6700 4200
rect 6900 4000 7000 4200
rect 5000 3600 5100 3800
rect 5300 3600 5400 3800
rect 5000 3500 5400 3600
rect 5425 3810 5535 3825
rect 5425 3790 5435 3810
rect 5455 3790 5505 3810
rect 5525 3790 5535 3810
rect 5425 3775 5535 3790
rect 5560 3810 6000 3825
rect 5560 3790 5570 3810
rect 5590 3790 6000 3810
rect 3395 3415 3405 3435
rect 3425 3415 3435 3435
rect 3395 3400 3435 3415
rect 3325 3270 3335 3290
rect 3355 3270 3365 3290
rect 3325 3260 3365 3270
rect 4500 3200 4900 3300
rect 4500 3000 4600 3200
rect 4800 3000 4900 3200
rect 4500 2900 4900 3000
rect 5100 2850 5300 3500
rect 5425 3290 5465 3775
rect 5495 3610 5535 3625
rect 5495 3590 5505 3610
rect 5525 3590 5535 3610
rect 5495 3435 5535 3590
rect 5560 3610 6000 3790
rect 5560 3590 5570 3610
rect 5590 3590 6000 3610
rect 5560 3575 6000 3590
rect 6600 3800 7000 4000
rect 6600 3600 6700 3800
rect 6900 3600 7000 3800
rect 6600 3500 7000 3600
rect 7100 3800 7500 4400
rect 7700 3825 8100 5300
rect 8200 5100 8600 5800
rect 8700 6000 9100 6200
rect 8700 5800 8800 6000
rect 9000 5800 9100 6000
rect 8700 5700 9100 5800
rect 10300 6000 10700 6100
rect 10300 5800 10400 6000
rect 10600 5800 10700 6000
rect 8700 5550 9100 5650
rect 8700 5350 8800 5550
rect 9000 5350 9100 5550
rect 8700 5250 9100 5350
rect 9800 5500 10200 5600
rect 9800 5300 9900 5500
rect 10100 5300 10200 5500
rect 8200 4900 8300 5100
rect 8500 4900 8600 5100
rect 8200 4200 8600 4900
rect 8700 5100 9100 5200
rect 8700 4900 8800 5100
rect 9000 4900 9100 5100
rect 8700 4650 9100 4900
rect 8700 4450 8800 4650
rect 9000 4450 9100 4650
rect 8700 4350 9100 4450
rect 9200 4600 9600 4700
rect 9200 4400 9300 4600
rect 9500 4400 9600 4600
rect 8200 4000 8300 4200
rect 8500 4000 8600 4200
rect 8200 3900 8600 4000
rect 8700 4200 9100 4300
rect 8700 4000 8800 4200
rect 9000 4000 9100 4200
rect 7100 3600 7200 3800
rect 7400 3600 7500 3800
rect 7100 3500 7500 3600
rect 7525 3810 7635 3825
rect 7525 3790 7535 3810
rect 7555 3790 7605 3810
rect 7625 3790 7635 3810
rect 7525 3775 7635 3790
rect 7660 3810 8100 3825
rect 7660 3790 7670 3810
rect 7690 3790 8100 3810
rect 5495 3415 5505 3435
rect 5525 3415 5535 3435
rect 5495 3400 5535 3415
rect 5425 3270 5435 3290
rect 5455 3270 5465 3290
rect 5425 3260 5465 3270
rect 6600 3200 7000 3300
rect 6600 3000 6700 3200
rect 6900 3000 7000 3200
rect 6600 2900 7000 3000
rect 7200 2850 7400 3500
rect 7525 3290 7565 3775
rect 7595 3610 7635 3625
rect 7595 3590 7605 3610
rect 7625 3590 7635 3610
rect 7595 3435 7635 3590
rect 7660 3610 8100 3790
rect 7660 3590 7670 3610
rect 7690 3590 8100 3610
rect 7660 3575 8100 3590
rect 8700 3800 9100 4000
rect 8700 3600 8800 3800
rect 9000 3600 9100 3800
rect 8700 3500 9100 3600
rect 9200 3800 9600 4400
rect 9800 3825 10200 5300
rect 10300 5100 10700 5800
rect 10900 6000 11300 6200
rect 10900 5800 11000 6000
rect 11200 5800 11300 6000
rect 10900 5700 11300 5800
rect 12500 6000 12900 6100
rect 12500 5800 12600 6000
rect 12800 5800 12900 6000
rect 10900 5550 11300 5650
rect 10900 5350 11000 5550
rect 11200 5350 11300 5550
rect 10900 5250 11300 5350
rect 12000 5500 12400 5600
rect 12000 5300 12100 5500
rect 12300 5300 12400 5500
rect 10300 4900 10400 5100
rect 10600 4900 10700 5100
rect 10300 4200 10700 4900
rect 10900 5100 11300 5200
rect 10900 4900 11000 5100
rect 11200 4900 11300 5100
rect 10900 4650 11300 4900
rect 10900 4450 11000 4650
rect 11200 4450 11300 4650
rect 10900 4350 11300 4450
rect 11400 4600 11800 4700
rect 11400 4400 11500 4600
rect 11700 4400 11800 4600
rect 10300 4000 10400 4200
rect 10600 4000 10700 4200
rect 10300 3900 10700 4000
rect 10900 4200 11300 4300
rect 10900 4000 11000 4200
rect 11200 4000 11300 4200
rect 9200 3600 9300 3800
rect 9500 3600 9600 3800
rect 9200 3500 9600 3600
rect 9625 3810 9735 3825
rect 9625 3790 9635 3810
rect 9655 3790 9705 3810
rect 9725 3790 9735 3810
rect 9625 3775 9735 3790
rect 9760 3810 10200 3825
rect 9760 3790 9770 3810
rect 9790 3790 10200 3810
rect 7595 3415 7605 3435
rect 7625 3415 7635 3435
rect 7595 3400 7635 3415
rect 7525 3270 7535 3290
rect 7555 3270 7565 3290
rect 7525 3260 7565 3270
rect 8700 3200 9100 3300
rect 8700 3000 8800 3200
rect 9000 3000 9100 3200
rect 8700 2900 9100 3000
rect 9300 2850 9500 3500
rect 9625 3290 9665 3775
rect 9695 3610 9735 3625
rect 9695 3590 9705 3610
rect 9725 3590 9735 3610
rect 9695 3435 9735 3590
rect 9760 3610 10200 3790
rect 9760 3590 9770 3610
rect 9790 3590 10200 3610
rect 9760 3575 10200 3590
rect 10900 3800 11300 4000
rect 10900 3600 11000 3800
rect 11200 3600 11300 3800
rect 10900 3500 11300 3600
rect 11400 3800 11800 4400
rect 12000 3825 12400 5300
rect 12500 5100 12900 5800
rect 13100 6000 13500 6200
rect 15600 6200 17100 6600
rect 13100 5800 13200 6000
rect 13400 5800 13500 6000
rect 13100 5700 13500 5800
rect 14700 6000 15100 6100
rect 14700 5800 14800 6000
rect 15000 5800 15100 6000
rect 13100 5550 13500 5650
rect 13100 5350 13200 5550
rect 13400 5350 13500 5550
rect 13100 5250 13500 5350
rect 14200 5500 14600 5600
rect 14200 5300 14300 5500
rect 14500 5300 14600 5500
rect 12500 4900 12600 5100
rect 12800 4900 12900 5100
rect 12500 4200 12900 4900
rect 13100 5100 13500 5200
rect 13100 4900 13200 5100
rect 13400 4900 13500 5100
rect 13100 4650 13500 4900
rect 13100 4450 13200 4650
rect 13400 4450 13500 4650
rect 13100 4350 13500 4450
rect 13600 4600 14000 4700
rect 13600 4400 13700 4600
rect 13900 4400 14000 4600
rect 12500 4000 12600 4200
rect 12800 4000 12900 4200
rect 12500 3900 12900 4000
rect 13100 4200 13500 4300
rect 13100 4000 13200 4200
rect 13400 4000 13500 4200
rect 11400 3600 11500 3800
rect 11700 3600 11800 3800
rect 11400 3500 11800 3600
rect 11825 3810 11935 3825
rect 11825 3790 11835 3810
rect 11855 3790 11905 3810
rect 11925 3790 11935 3810
rect 11825 3775 11935 3790
rect 11960 3810 12400 3825
rect 11960 3790 11970 3810
rect 11990 3790 12400 3810
rect 9695 3415 9705 3435
rect 9725 3415 9735 3435
rect 9695 3400 9735 3415
rect 9625 3270 9635 3290
rect 9655 3270 9665 3290
rect 9625 3260 9665 3270
rect 10900 3200 11300 3300
rect 10900 3000 11000 3200
rect 11200 3000 11300 3200
rect 10900 2900 11300 3000
rect 11500 2850 11700 3500
rect 11825 3290 11865 3775
rect 11895 3610 11935 3625
rect 11895 3590 11905 3610
rect 11925 3590 11935 3610
rect 11895 3435 11935 3590
rect 11960 3610 12400 3790
rect 11960 3590 11970 3610
rect 11990 3590 12400 3610
rect 11960 3575 12400 3590
rect 13100 3800 13500 4000
rect 13100 3600 13200 3800
rect 13400 3600 13500 3800
rect 13100 3500 13500 3600
rect 13600 3800 14000 4400
rect 14200 3825 14600 5300
rect 14700 5100 15100 5800
rect 15150 5550 15550 5650
rect 15150 5350 15250 5550
rect 15450 5350 15550 5550
rect 15150 5250 15550 5350
rect 14700 4900 14800 5100
rect 15000 4900 15100 5100
rect 14700 4200 15100 4900
rect 14700 4000 14800 4200
rect 15000 4000 15100 4200
rect 14700 3900 15100 4000
rect 13600 3600 13700 3800
rect 13900 3600 14000 3800
rect 13600 3500 14000 3600
rect 14025 3810 14135 3825
rect 14025 3790 14035 3810
rect 14055 3790 14105 3810
rect 14125 3790 14135 3810
rect 14025 3775 14135 3790
rect 14160 3810 14600 3825
rect 14160 3790 14170 3810
rect 14190 3790 14600 3810
rect 11895 3415 11905 3435
rect 11925 3415 11935 3435
rect 11895 3400 11935 3415
rect 11825 3270 11835 3290
rect 11855 3270 11865 3290
rect 11825 3260 11865 3270
rect 13100 3200 13500 3300
rect 13100 3000 13200 3200
rect 13400 3000 13500 3200
rect 13100 2900 13500 3000
rect 13700 2850 13900 3500
rect 14025 3290 14065 3775
rect 14095 3610 14135 3625
rect 14095 3590 14105 3610
rect 14125 3590 14135 3610
rect 14095 3435 14135 3590
rect 14160 3610 14600 3790
rect 14160 3590 14170 3610
rect 14190 3590 14600 3610
rect 14160 3575 14600 3590
rect 15600 3800 16000 6200
rect 15600 3600 15700 3800
rect 15900 3600 16000 3800
rect 15600 3500 16000 3600
rect 14095 3415 14105 3435
rect 14125 3415 14135 3435
rect 14095 3400 14135 3415
rect 14025 3270 14035 3290
rect 14055 3270 14065 3290
rect 14025 3260 14065 3270
rect 15150 3200 15550 3300
rect 15150 3000 15250 3200
rect 15450 3000 15550 3200
rect 15150 2900 15550 3000
<< viali >>
rect 400 7750 600 7950
rect 2300 7750 2500 7950
rect 4400 7750 4600 7950
rect 6500 7750 6700 7950
rect 8600 7750 8800 7950
rect 10700 7750 10900 7950
rect 12900 7750 13100 7950
rect 15000 7750 15200 7950
rect 16800 7750 17000 7950
rect 400 5350 600 5550
rect 400 4450 600 4650
rect 400 3600 600 3800
rect 2500 5350 2700 5550
rect 2500 4450 2700 4650
rect 400 3000 600 3200
rect 2500 3600 2700 3800
rect 4600 5350 4800 5550
rect 4600 4450 4800 4650
rect 1305 3415 1325 3435
rect 1235 3270 1255 3290
rect 2500 3000 2700 3200
rect 4600 3600 4800 3800
rect 6700 5350 6900 5550
rect 6700 4450 6900 4650
rect 3405 3415 3425 3435
rect 3335 3270 3355 3290
rect 4600 3000 4800 3200
rect 6700 3600 6900 3800
rect 8800 5350 9000 5550
rect 8800 4450 9000 4650
rect 5505 3415 5525 3435
rect 5435 3270 5455 3290
rect 6700 3000 6900 3200
rect 8800 3600 9000 3800
rect 11000 5350 11200 5550
rect 11000 4450 11200 4650
rect 7605 3415 7625 3435
rect 7535 3270 7555 3290
rect 8800 3000 9000 3200
rect 11000 3600 11200 3800
rect 13200 5350 13400 5550
rect 13200 4450 13400 4650
rect 9705 3415 9725 3435
rect 9635 3270 9655 3290
rect 11000 3000 11200 3200
rect 13200 3600 13400 3800
rect 15250 5350 15450 5550
rect 11905 3415 11925 3435
rect 11835 3270 11855 3290
rect 13200 3000 13400 3200
rect 15700 3600 15900 3800
rect 14105 3415 14125 3435
rect 14035 3270 14055 3290
rect 15250 3000 15450 3200
<< metal1 >>
rect 300 7950 17550 8050
rect 300 7750 400 7950
rect 600 7750 2300 7950
rect 2500 7750 4400 7950
rect 4600 7750 6500 7950
rect 6700 7750 8600 7950
rect 8800 7750 10700 7950
rect 10900 7750 12900 7950
rect 13100 7750 15000 7950
rect 15200 7750 16800 7950
rect 17000 7750 17550 7950
rect 300 7650 17550 7750
rect 17150 5650 17550 7650
rect -100 5550 17550 5650
rect -100 5350 400 5550
rect 600 5350 2500 5550
rect 2700 5350 4600 5550
rect 4800 5350 6700 5550
rect 6900 5350 8800 5550
rect 9000 5350 11000 5550
rect 11200 5350 13200 5550
rect 13400 5350 15250 5550
rect 15450 5350 17550 5550
rect -100 5250 17550 5350
rect -100 3300 250 5250
rect 300 4650 16000 4750
rect 300 4450 400 4650
rect 600 4600 2500 4650
rect 600 4450 900 4600
rect 300 4400 900 4450
rect 1100 4450 2500 4600
rect 2700 4450 4600 4650
rect 4800 4450 6700 4650
rect 6900 4450 8800 4650
rect 9000 4450 11000 4650
rect 11200 4450 13200 4650
rect 13400 4450 16000 4650
rect 1100 4400 16000 4450
rect 300 4350 16000 4400
rect 300 3800 16000 3900
rect 300 3600 400 3800
rect 600 3600 2500 3800
rect 2700 3600 4600 3800
rect 4800 3600 6700 3800
rect 6900 3600 8800 3800
rect 9000 3600 11000 3800
rect 11200 3600 13200 3800
rect 13400 3600 15700 3800
rect 15900 3600 16000 3800
rect 300 3500 16000 3600
rect 300 3435 16000 3450
rect 300 3415 1305 3435
rect 1325 3415 3405 3435
rect 3425 3415 5505 3435
rect 5525 3415 7605 3435
rect 7625 3415 9705 3435
rect 9725 3415 11905 3435
rect 11925 3415 14105 3435
rect 14125 3415 16000 3435
rect 300 3350 16000 3415
rect -100 3290 15550 3300
rect -100 3270 1235 3290
rect 1255 3270 3335 3290
rect 3355 3270 5435 3290
rect 5455 3270 7535 3290
rect 7555 3270 9635 3290
rect 9655 3270 11835 3290
rect 11855 3270 14035 3290
rect 14055 3270 15550 3290
rect -100 3200 15550 3270
rect -100 3000 400 3200
rect 600 3000 2500 3200
rect 2700 3000 4600 3200
rect 4800 3000 6700 3200
rect 6900 3000 8800 3200
rect 9000 3000 11000 3200
rect 11200 3000 13200 3200
rect 13400 3000 15250 3200
rect 15450 3000 15550 3200
rect -100 2900 15550 3000
<< labels >>
rlabel metal1 -100 2900 -100 5650 7 VP
port 4 w
rlabel locali -50 6200 -50 6600 7 IIN
port 6 w
rlabel poly -100 6200 -100 6600 7 VGATE
port 13 w
rlabel locali 3000 2850 3200 2850 5 D5
port 7 s
rlabel locali 5100 2850 5300 2850 5 D4
port 8 s
rlabel locali 7200 2850 7400 2850 5 D3
port 9 s
rlabel locali 9300 2850 9500 2850 5 D2
port 10 s
rlabel locali 11500 2850 11700 2850 5 D1
port 11 s
rlabel metal1 16000 3350 16000 3450 3 VN
port 2 e
rlabel locali 13700 2850 13900 2850 5 D0
port 12 s
rlabel locali 900 2850 1100 2850 5 D6
port 5 s
rlabel metal1 16000 3500 16000 3900 3 IDUMP
port 14 e
rlabel metal1 16000 4350 16000 4750 3 IOUT
port 15 e
<< end >>
