magic
tech sky130A
timestamp 1763024294
<< nwell >>
rect -1000 -700 33950 2400
<< pmos >>
rect 0 1900 1200 2300
rect 2500 1900 3700 2300
rect 5000 1900 6200 2300
rect 7500 1900 8700 2300
rect 10000 1900 11200 2300
rect 12500 1900 13700 2300
rect 15000 1900 16200 2300
rect 17500 1900 18700 2300
rect 20000 1900 21200 2300
rect 22500 1900 23700 2300
rect 25000 1900 26200 2300
rect 27500 1900 28700 2300
rect 30000 1900 31200 2300
rect 0 1400 1200 1800
rect 2500 1400 3700 1800
rect 5000 1400 6200 1800
rect 7500 1400 8700 1800
rect 10000 1400 11200 1800
rect 12500 1400 13700 1800
rect 15000 1400 16200 1800
rect 17500 1400 18700 1800
rect 20000 1400 21200 1800
rect 22500 1400 23700 1800
rect 25000 1400 26200 1800
rect 27500 1400 28700 1800
rect 30000 1400 31200 1800
rect 32000 1400 33200 1800
rect 0 900 1200 1300
rect 2500 900 3700 1300
rect 5000 900 6200 1300
rect 7500 900 8700 1300
rect 10000 900 11200 1300
rect 12500 900 13700 1300
rect 15000 900 16200 1300
rect 17500 900 18700 1300
rect 20000 900 21200 1300
rect 22500 900 23700 1300
rect 25000 900 26200 1300
rect 27500 900 28700 1300
rect 30000 900 31200 1300
rect 32000 900 33200 1300
rect 0 -100 1200 300
rect 2500 -100 3700 300
rect 5000 -100 6200 300
rect 7500 -100 8700 300
rect 10000 -100 11200 300
rect 12500 -100 13700 300
rect 15000 -100 16200 300
rect 17500 -100 18700 300
rect 20000 -100 21200 300
rect 22500 -100 23700 300
rect 25000 -100 26200 300
rect 27500 -100 28700 300
rect 30000 -100 31200 300
rect 0 -600 1200 -200
rect 2500 -600 3700 -200
rect 5000 -600 6200 -200
rect 7500 -600 8700 -200
rect 10000 -600 11200 -200
rect 12500 -600 13700 -200
rect 15000 -600 16200 -200
rect 17500 -600 18700 -200
rect 20000 -600 21200 -200
rect 22500 -600 23700 -200
rect 25000 -600 26200 -200
rect 27500 -600 28700 -200
rect 30000 -600 31200 -200
<< pdiff >>
rect -400 2200 0 2300
rect -400 2000 -300 2200
rect -100 2000 0 2200
rect -400 1900 0 2000
rect 1200 2200 1600 2300
rect 2100 2200 2500 2300
rect 1200 2000 1300 2200
rect 1500 2000 1600 2200
rect 2100 2000 2200 2200
rect 2400 2000 2500 2200
rect 1200 1900 1600 2000
rect 2100 1900 2500 2000
rect 3700 2200 4100 2300
rect 4600 2200 5000 2300
rect 3700 2000 3800 2200
rect 4000 2000 4100 2200
rect 4600 2000 4700 2200
rect 4900 2000 5000 2200
rect 3700 1900 4100 2000
rect 4600 1900 5000 2000
rect 6200 2200 6600 2300
rect 7100 2200 7500 2300
rect 6200 2000 6300 2200
rect 6500 2000 6600 2200
rect 7100 2000 7200 2200
rect 7400 2000 7500 2200
rect 6200 1900 6600 2000
rect 7100 1900 7500 2000
rect 8700 2200 9100 2300
rect 9600 2200 10000 2300
rect 8700 2000 8800 2200
rect 9000 2000 9100 2200
rect 9600 2000 9700 2200
rect 9900 2000 10000 2200
rect 8700 1900 9100 2000
rect 9600 1900 10000 2000
rect 11200 2200 11600 2300
rect 12100 2200 12500 2300
rect 11200 2000 11300 2200
rect 11500 2000 11600 2200
rect 12100 2000 12200 2200
rect 12400 2000 12500 2200
rect 11200 1900 11600 2000
rect 12100 1900 12500 2000
rect 13700 2200 14100 2300
rect 14600 2200 15000 2300
rect 13700 2000 13800 2200
rect 14000 2000 14100 2200
rect 14600 2000 14700 2200
rect 14900 2000 15000 2200
rect 13700 1900 14100 2000
rect 14600 1900 15000 2000
rect 16200 2200 16600 2300
rect 17100 2200 17500 2300
rect 16200 2000 16300 2200
rect 16500 2000 16600 2200
rect 17100 2000 17200 2200
rect 17400 2000 17500 2200
rect 16200 1900 16600 2000
rect 17100 1900 17500 2000
rect 18700 2200 19100 2300
rect 19600 2200 20000 2300
rect 18700 2000 18800 2200
rect 19000 2000 19100 2200
rect 19600 2000 19700 2200
rect 19900 2000 20000 2200
rect 18700 1900 19100 2000
rect 19600 1900 20000 2000
rect 21200 2200 21600 2300
rect 22100 2200 22500 2300
rect 21200 2000 21300 2200
rect 21500 2000 21600 2200
rect 22100 2000 22200 2200
rect 22400 2000 22500 2200
rect 21200 1900 21600 2000
rect 22100 1900 22500 2000
rect 23700 2200 24100 2300
rect 24600 2200 25000 2300
rect 23700 2000 23800 2200
rect 24000 2000 24100 2200
rect 24600 2000 24700 2200
rect 24900 2000 25000 2200
rect 23700 1900 24100 2000
rect 24600 1900 25000 2000
rect 26200 2200 26600 2300
rect 27100 2200 27500 2300
rect 26200 2000 26300 2200
rect 26500 2000 26600 2200
rect 27100 2000 27200 2200
rect 27400 2000 27500 2200
rect 26200 1900 26600 2000
rect 27100 1900 27500 2000
rect 28700 2200 29100 2300
rect 29600 2200 30000 2300
rect 28700 2000 28800 2200
rect 29000 2000 29100 2200
rect 29600 2000 29700 2200
rect 29900 2000 30000 2200
rect 28700 1900 29100 2000
rect 29600 1900 30000 2000
rect 31200 2200 31600 2300
rect 31200 2000 31300 2200
rect 31500 2000 31600 2200
rect 31200 1900 31600 2000
rect -400 1700 0 1800
rect -400 1500 -300 1700
rect -100 1500 0 1700
rect -400 1400 0 1500
rect 1200 1700 1600 1800
rect 1200 1500 1300 1700
rect 1500 1500 1600 1700
rect 1200 1400 1600 1500
rect 2100 1700 2500 1800
rect 2100 1500 2200 1700
rect 2400 1500 2500 1700
rect 2100 1400 2500 1500
rect 3700 1700 4100 1800
rect 3700 1500 3800 1700
rect 4000 1500 4100 1700
rect 3700 1400 4100 1500
rect 4600 1700 5000 1800
rect 4600 1500 4700 1700
rect 4900 1500 5000 1700
rect 4600 1400 5000 1500
rect 6200 1700 6600 1800
rect 6200 1500 6300 1700
rect 6500 1500 6600 1700
rect 6200 1400 6600 1500
rect 7100 1700 7500 1800
rect 7100 1500 7200 1700
rect 7400 1500 7500 1700
rect 7100 1400 7500 1500
rect 8700 1700 9100 1800
rect 8700 1500 8800 1700
rect 9000 1500 9100 1700
rect 8700 1400 9100 1500
rect 9600 1700 10000 1800
rect 9600 1500 9700 1700
rect 9900 1500 10000 1700
rect 9600 1400 10000 1500
rect 11200 1700 11600 1800
rect 11200 1500 11300 1700
rect 11500 1500 11600 1700
rect 11200 1400 11600 1500
rect 12100 1700 12500 1800
rect 12100 1500 12200 1700
rect 12400 1500 12500 1700
rect 12100 1400 12500 1500
rect 13700 1700 14100 1800
rect 13700 1500 13800 1700
rect 14000 1500 14100 1700
rect 13700 1400 14100 1500
rect 14600 1700 15000 1800
rect 14600 1500 14700 1700
rect 14900 1500 15000 1700
rect 14600 1400 15000 1500
rect 16200 1700 16600 1800
rect 16200 1500 16300 1700
rect 16500 1500 16600 1700
rect 16200 1400 16600 1500
rect 17100 1700 17500 1800
rect 17100 1500 17200 1700
rect 17400 1500 17500 1700
rect 17100 1400 17500 1500
rect 18700 1700 19100 1800
rect 18700 1500 18800 1700
rect 19000 1500 19100 1700
rect 18700 1400 19100 1500
rect 19600 1700 20000 1800
rect 19600 1500 19700 1700
rect 19900 1500 20000 1700
rect 19600 1400 20000 1500
rect 21200 1700 21600 1800
rect 21200 1500 21300 1700
rect 21500 1500 21600 1700
rect 21200 1400 21600 1500
rect 22100 1700 22500 1800
rect 22100 1500 22200 1700
rect 22400 1500 22500 1700
rect 22100 1400 22500 1500
rect 23700 1700 24100 1800
rect 23700 1500 23800 1700
rect 24000 1500 24100 1700
rect 23700 1400 24100 1500
rect 24600 1700 25000 1800
rect 24600 1500 24700 1700
rect 24900 1500 25000 1700
rect 24600 1400 25000 1500
rect 26200 1700 26600 1800
rect 26200 1500 26300 1700
rect 26500 1500 26600 1700
rect 26200 1400 26600 1500
rect 27100 1700 27500 1800
rect 27100 1500 27200 1700
rect 27400 1500 27500 1700
rect 27100 1400 27500 1500
rect 28700 1700 29100 1800
rect 28700 1500 28800 1700
rect 29000 1500 29100 1700
rect 28700 1400 29100 1500
rect 29600 1700 30000 1800
rect 29600 1500 29700 1700
rect 29900 1500 30000 1700
rect 29600 1400 30000 1500
rect 31200 1700 32000 1800
rect 31200 1500 31300 1700
rect 31500 1500 31700 1700
rect 31900 1500 32000 1700
rect 31200 1400 32000 1500
rect 33200 1700 33600 1800
rect 33200 1500 33300 1700
rect 33500 1500 33600 1700
rect 33200 1400 33600 1500
rect -400 1200 0 1300
rect -400 1000 -300 1200
rect -100 1000 0 1200
rect -400 900 0 1000
rect 1200 1200 1600 1300
rect 1200 1000 1300 1200
rect 1500 1000 1600 1200
rect 1200 900 1600 1000
rect 2100 1200 2500 1300
rect 2100 1000 2200 1200
rect 2400 1000 2500 1200
rect 2100 900 2500 1000
rect 3700 1200 4100 1300
rect 3700 1000 3800 1200
rect 4000 1000 4100 1200
rect 3700 900 4100 1000
rect 4600 1200 5000 1300
rect 4600 1000 4700 1200
rect 4900 1000 5000 1200
rect 4600 900 5000 1000
rect 6200 1200 6600 1300
rect 6200 1000 6300 1200
rect 6500 1000 6600 1200
rect 6200 900 6600 1000
rect 7100 1200 7500 1300
rect 7100 1000 7200 1200
rect 7400 1000 7500 1200
rect 7100 900 7500 1000
rect 8700 1200 9100 1300
rect 8700 1000 8800 1200
rect 9000 1000 9100 1200
rect 8700 900 9100 1000
rect 9600 1200 10000 1300
rect 9600 1000 9700 1200
rect 9900 1000 10000 1200
rect 9600 900 10000 1000
rect 11200 1200 11600 1300
rect 11200 1000 11300 1200
rect 11500 1000 11600 1200
rect 11200 900 11600 1000
rect 12100 1200 12500 1300
rect 12100 1000 12200 1200
rect 12400 1000 12500 1200
rect 12100 900 12500 1000
rect 13700 1200 14100 1300
rect 13700 1000 13800 1200
rect 14000 1000 14100 1200
rect 13700 900 14100 1000
rect 14600 1200 15000 1300
rect 14600 1000 14700 1200
rect 14900 1000 15000 1200
rect 14600 900 15000 1000
rect 16200 1200 16600 1300
rect 16200 1000 16300 1200
rect 16500 1000 16600 1200
rect 16200 900 16600 1000
rect 17100 1200 17500 1300
rect 17100 1000 17200 1200
rect 17400 1000 17500 1200
rect 17100 900 17500 1000
rect 18700 1200 19100 1300
rect 18700 1000 18800 1200
rect 19000 1000 19100 1200
rect 18700 900 19100 1000
rect 19600 1200 20000 1300
rect 19600 1000 19700 1200
rect 19900 1000 20000 1200
rect 19600 900 20000 1000
rect 21200 1200 21600 1300
rect 21200 1000 21300 1200
rect 21500 1000 21600 1200
rect 21200 900 21600 1000
rect 22100 1200 22500 1300
rect 22100 1000 22200 1200
rect 22400 1000 22500 1200
rect 22100 900 22500 1000
rect 23700 1200 24100 1300
rect 23700 1000 23800 1200
rect 24000 1000 24100 1200
rect 23700 900 24100 1000
rect 24600 1200 25000 1300
rect 24600 1000 24700 1200
rect 24900 1000 25000 1200
rect 24600 900 25000 1000
rect 26200 1200 26600 1300
rect 26200 1000 26300 1200
rect 26500 1000 26600 1200
rect 26200 900 26600 1000
rect 27100 1200 27500 1300
rect 27100 1000 27200 1200
rect 27400 1000 27500 1200
rect 27100 900 27500 1000
rect 28700 1200 29100 1300
rect 28700 1000 28800 1200
rect 29000 1000 29100 1200
rect 28700 900 29100 1000
rect 29600 1200 30000 1300
rect 29600 1000 29700 1200
rect 29900 1000 30000 1200
rect 29600 900 30000 1000
rect 31200 1200 32000 1300
rect 31200 1000 31300 1200
rect 31500 1000 31700 1200
rect 31900 1000 32000 1200
rect 31200 900 32000 1000
rect 33200 1200 33600 1300
rect 33200 1000 33300 1200
rect 33500 1000 33600 1200
rect 33200 900 33600 1000
rect -400 200 0 300
rect -400 0 -300 200
rect -100 0 0 200
rect -400 -100 0 0
rect 1200 200 1600 300
rect 1200 0 1300 200
rect 1500 0 1600 200
rect 1200 -100 1600 0
rect 2100 200 2500 300
rect 2100 0 2200 200
rect 2400 0 2500 200
rect 2100 -100 2500 0
rect 3700 200 4100 300
rect 3700 0 3800 200
rect 4000 0 4100 200
rect 3700 -100 4100 0
rect 4600 200 5000 300
rect 4600 0 4700 200
rect 4900 0 5000 200
rect 4600 -100 5000 0
rect 6200 200 6600 300
rect 6200 0 6300 200
rect 6500 0 6600 200
rect 6200 -100 6600 0
rect 7100 200 7500 300
rect 7100 0 7200 200
rect 7400 0 7500 200
rect 7100 -100 7500 0
rect 8700 200 9100 300
rect 8700 0 8800 200
rect 9000 0 9100 200
rect 8700 -100 9100 0
rect 9600 200 10000 300
rect 9600 0 9700 200
rect 9900 0 10000 200
rect 9600 -100 10000 0
rect 11200 200 11600 300
rect 11200 0 11300 200
rect 11500 0 11600 200
rect 11200 -100 11600 0
rect 12100 200 12500 300
rect 12100 0 12200 200
rect 12400 0 12500 200
rect 12100 -100 12500 0
rect 13700 200 14100 300
rect 13700 0 13800 200
rect 14000 0 14100 200
rect 13700 -100 14100 0
rect 14600 200 15000 300
rect 14600 0 14700 200
rect 14900 0 15000 200
rect 14600 -100 15000 0
rect 16200 200 16600 300
rect 16200 0 16300 200
rect 16500 0 16600 200
rect 16200 -100 16600 0
rect 17100 200 17500 300
rect 17100 0 17200 200
rect 17400 0 17500 200
rect 17100 -100 17500 0
rect 18700 200 19100 300
rect 18700 0 18800 200
rect 19000 0 19100 200
rect 18700 -100 19100 0
rect 19600 200 20000 300
rect 19600 0 19700 200
rect 19900 0 20000 200
rect 19600 -100 20000 0
rect 21200 200 21600 300
rect 21200 0 21300 200
rect 21500 0 21600 200
rect 21200 -100 21600 0
rect 22100 200 22500 300
rect 22100 0 22200 200
rect 22400 0 22500 200
rect 22100 -100 22500 0
rect 23700 200 24100 300
rect 23700 0 23800 200
rect 24000 0 24100 200
rect 23700 -100 24100 0
rect 24600 200 25000 300
rect 24600 0 24700 200
rect 24900 0 25000 200
rect 24600 -100 25000 0
rect 26200 200 26600 300
rect 26200 0 26300 200
rect 26500 0 26600 200
rect 26200 -100 26600 0
rect 27100 200 27500 300
rect 27100 0 27200 200
rect 27400 0 27500 200
rect 27100 -100 27500 0
rect 28700 200 29100 300
rect 28700 0 28800 200
rect 29000 0 29100 200
rect 28700 -100 29100 0
rect 29600 200 30000 300
rect 29600 0 29700 200
rect 29900 0 30000 200
rect 29600 -100 30000 0
rect 31200 200 31600 300
rect 31200 0 31300 200
rect 31500 0 31600 200
rect 31200 -100 31600 0
rect -400 -300 0 -200
rect -400 -500 -300 -300
rect -100 -500 0 -300
rect -400 -600 0 -500
rect 1200 -300 1600 -200
rect 2100 -300 2500 -200
rect 1200 -500 1300 -300
rect 1500 -500 1600 -300
rect 2100 -500 2200 -300
rect 2400 -500 2500 -300
rect 1200 -600 1600 -500
rect 2100 -600 2500 -500
rect 3700 -300 4100 -200
rect 4600 -300 5000 -200
rect 3700 -500 3800 -300
rect 4000 -500 4100 -300
rect 4600 -500 4700 -300
rect 4900 -500 5000 -300
rect 3700 -600 4100 -500
rect 4600 -600 5000 -500
rect 6200 -300 6600 -200
rect 7100 -300 7500 -200
rect 6200 -500 6300 -300
rect 6500 -500 6600 -300
rect 7100 -500 7200 -300
rect 7400 -500 7500 -300
rect 6200 -600 6600 -500
rect 7100 -600 7500 -500
rect 8700 -300 9100 -200
rect 9600 -300 10000 -200
rect 8700 -500 8800 -300
rect 9000 -500 9100 -300
rect 9600 -500 9700 -300
rect 9900 -500 10000 -300
rect 8700 -600 9100 -500
rect 9600 -600 10000 -500
rect 11200 -300 11600 -200
rect 12100 -300 12500 -200
rect 11200 -500 11300 -300
rect 11500 -500 11600 -300
rect 12100 -500 12200 -300
rect 12400 -500 12500 -300
rect 11200 -600 11600 -500
rect 12100 -600 12500 -500
rect 13700 -300 14100 -200
rect 14600 -300 15000 -200
rect 13700 -500 13800 -300
rect 14000 -500 14100 -300
rect 14600 -500 14700 -300
rect 14900 -500 15000 -300
rect 13700 -600 14100 -500
rect 14600 -600 15000 -500
rect 16200 -300 16600 -200
rect 17100 -300 17500 -200
rect 16200 -500 16300 -300
rect 16500 -500 16600 -300
rect 17100 -500 17200 -300
rect 17400 -500 17500 -300
rect 16200 -600 16600 -500
rect 17100 -600 17500 -500
rect 18700 -300 19100 -200
rect 19600 -300 20000 -200
rect 18700 -500 18800 -300
rect 19000 -500 19100 -300
rect 19600 -500 19700 -300
rect 19900 -500 20000 -300
rect 18700 -600 19100 -500
rect 19600 -600 20000 -500
rect 21200 -300 21600 -200
rect 22100 -300 22500 -200
rect 21200 -500 21300 -300
rect 21500 -500 21600 -300
rect 22100 -500 22200 -300
rect 22400 -500 22500 -300
rect 21200 -600 21600 -500
rect 22100 -600 22500 -500
rect 23700 -300 24100 -200
rect 24600 -300 25000 -200
rect 23700 -500 23800 -300
rect 24000 -500 24100 -300
rect 24600 -500 24700 -300
rect 24900 -500 25000 -300
rect 23700 -600 24100 -500
rect 24600 -600 25000 -500
rect 26200 -300 26600 -200
rect 27100 -300 27500 -200
rect 26200 -500 26300 -300
rect 26500 -500 26600 -300
rect 27100 -500 27200 -300
rect 27400 -500 27500 -300
rect 26200 -600 26600 -500
rect 27100 -600 27500 -500
rect 28700 -300 29100 -200
rect 29600 -300 30000 -200
rect 28700 -500 28800 -300
rect 29000 -500 29100 -300
rect 29600 -500 29700 -300
rect 29900 -500 30000 -300
rect 28700 -600 29100 -500
rect 29600 -600 30000 -500
rect 31200 -300 31600 -200
rect 31200 -500 31300 -300
rect 31500 -500 31600 -300
rect 31200 -600 31600 -500
<< pdiffc >>
rect -300 2000 -100 2200
rect 1300 2000 1500 2200
rect 2200 2000 2400 2200
rect 3800 2000 4000 2200
rect 4700 2000 4900 2200
rect 6300 2000 6500 2200
rect 7200 2000 7400 2200
rect 8800 2000 9000 2200
rect 9700 2000 9900 2200
rect 11300 2000 11500 2200
rect 12200 2000 12400 2200
rect 13800 2000 14000 2200
rect 14700 2000 14900 2200
rect 16300 2000 16500 2200
rect 17200 2000 17400 2200
rect 18800 2000 19000 2200
rect 19700 2000 19900 2200
rect 21300 2000 21500 2200
rect 22200 2000 22400 2200
rect 23800 2000 24000 2200
rect 24700 2000 24900 2200
rect 26300 2000 26500 2200
rect 27200 2000 27400 2200
rect 28800 2000 29000 2200
rect 29700 2000 29900 2200
rect 31300 2000 31500 2200
rect -300 1500 -100 1700
rect 1300 1500 1500 1700
rect 2200 1500 2400 1700
rect 3800 1500 4000 1700
rect 4700 1500 4900 1700
rect 6300 1500 6500 1700
rect 7200 1500 7400 1700
rect 8800 1500 9000 1700
rect 9700 1500 9900 1700
rect 11300 1500 11500 1700
rect 12200 1500 12400 1700
rect 13800 1500 14000 1700
rect 14700 1500 14900 1700
rect 16300 1500 16500 1700
rect 17200 1500 17400 1700
rect 18800 1500 19000 1700
rect 19700 1500 19900 1700
rect 21300 1500 21500 1700
rect 22200 1500 22400 1700
rect 23800 1500 24000 1700
rect 24700 1500 24900 1700
rect 26300 1500 26500 1700
rect 27200 1500 27400 1700
rect 28800 1500 29000 1700
rect 29700 1500 29900 1700
rect 31300 1500 31500 1700
rect 31700 1500 31900 1700
rect 33300 1500 33500 1700
rect -300 1000 -100 1200
rect 1300 1000 1500 1200
rect 2200 1000 2400 1200
rect 3800 1000 4000 1200
rect 4700 1000 4900 1200
rect 6300 1000 6500 1200
rect 7200 1000 7400 1200
rect 8800 1000 9000 1200
rect 9700 1000 9900 1200
rect 11300 1000 11500 1200
rect 12200 1000 12400 1200
rect 13800 1000 14000 1200
rect 14700 1000 14900 1200
rect 16300 1000 16500 1200
rect 17200 1000 17400 1200
rect 18800 1000 19000 1200
rect 19700 1000 19900 1200
rect 21300 1000 21500 1200
rect 22200 1000 22400 1200
rect 23800 1000 24000 1200
rect 24700 1000 24900 1200
rect 26300 1000 26500 1200
rect 27200 1000 27400 1200
rect 28800 1000 29000 1200
rect 29700 1000 29900 1200
rect 31300 1000 31500 1200
rect 31700 1000 31900 1200
rect 33300 1000 33500 1200
rect -300 0 -100 200
rect 1300 0 1500 200
rect 2200 0 2400 200
rect 3800 0 4000 200
rect 4700 0 4900 200
rect 6300 0 6500 200
rect 7200 0 7400 200
rect 8800 0 9000 200
rect 9700 0 9900 200
rect 11300 0 11500 200
rect 12200 0 12400 200
rect 13800 0 14000 200
rect 14700 0 14900 200
rect 16300 0 16500 200
rect 17200 0 17400 200
rect 18800 0 19000 200
rect 19700 0 19900 200
rect 21300 0 21500 200
rect 22200 0 22400 200
rect 23800 0 24000 200
rect 24700 0 24900 200
rect 26300 0 26500 200
rect 27200 0 27400 200
rect 28800 0 29000 200
rect 29700 0 29900 200
rect 31300 0 31500 200
rect -300 -500 -100 -300
rect 1300 -500 1500 -300
rect 2200 -500 2400 -300
rect 3800 -500 4000 -300
rect 4700 -500 4900 -300
rect 6300 -500 6500 -300
rect 7200 -500 7400 -300
rect 8800 -500 9000 -300
rect 9700 -500 9900 -300
rect 11300 -500 11500 -300
rect 12200 -500 12400 -300
rect 13800 -500 14000 -300
rect 14700 -500 14900 -300
rect 16300 -500 16500 -300
rect 17200 -500 17400 -300
rect 18800 -500 19000 -300
rect 19700 -500 19900 -300
rect 21300 -500 21500 -300
rect 22200 -500 22400 -300
rect 23800 -500 24000 -300
rect 24700 -500 24900 -300
rect 26300 -500 26500 -300
rect 27200 -500 27400 -300
rect 28800 -500 29000 -300
rect 29700 -500 29900 -300
rect 31300 -500 31500 -300
<< nsubdiff >>
rect -900 2200 -400 2300
rect -900 2000 -800 2200
rect -600 2000 -400 2200
rect -900 1900 -400 2000
rect 1600 2200 2100 2300
rect 1600 2000 1750 2200
rect 1950 2000 2100 2200
rect 1600 1900 2100 2000
rect 4100 2200 4600 2300
rect 4100 2000 4250 2200
rect 4450 2000 4600 2200
rect 4100 1900 4600 2000
rect 6600 2200 7100 2300
rect 6600 2000 6750 2200
rect 6950 2000 7100 2200
rect 6600 1900 7100 2000
rect 9100 2200 9600 2300
rect 9100 2000 9250 2200
rect 9450 2000 9600 2200
rect 9100 1900 9600 2000
rect 11600 2200 12100 2300
rect 11600 2000 11750 2200
rect 11950 2000 12100 2200
rect 11600 1900 12100 2000
rect 14100 2200 14600 2300
rect 14100 2000 14250 2200
rect 14450 2000 14600 2200
rect 14100 1900 14600 2000
rect 16600 2200 17100 2300
rect 16600 2000 16750 2200
rect 16950 2000 17100 2200
rect 16600 1900 17100 2000
rect 19100 2200 19600 2300
rect 19100 2000 19250 2200
rect 19450 2000 19600 2200
rect 19100 1900 19600 2000
rect 21600 2200 22100 2300
rect 21600 2000 21750 2200
rect 21950 2000 22100 2200
rect 21600 1900 22100 2000
rect 24100 2200 24600 2300
rect 24100 2000 24250 2200
rect 24450 2000 24600 2200
rect 24100 1900 24600 2000
rect 26600 2200 27100 2300
rect 26600 2000 26750 2200
rect 26950 2000 27100 2200
rect 26600 1900 27100 2000
rect 29100 2200 29600 2300
rect 29100 2000 29250 2200
rect 29450 2000 29600 2200
rect 29100 1900 29600 2000
rect 31600 2200 32000 2300
rect 31600 2000 31700 2200
rect 31900 2000 32000 2200
rect 31600 1900 32000 2000
rect 33200 2200 33600 2300
rect 33200 2000 33300 2200
rect 33500 2000 33600 2200
rect 33200 1900 33600 2000
rect -900 -300 -400 -200
rect -900 -500 -800 -300
rect -600 -500 -400 -300
rect -900 -600 -400 -500
rect 1600 -300 2100 -200
rect 1600 -500 1750 -300
rect 1950 -500 2100 -300
rect 1600 -600 2100 -500
rect 4100 -300 4600 -200
rect 4100 -500 4250 -300
rect 4450 -500 4600 -300
rect 4100 -600 4600 -500
rect 6600 -300 7100 -200
rect 6600 -500 6750 -300
rect 6950 -500 7100 -300
rect 6600 -600 7100 -500
rect 9100 -300 9600 -200
rect 9100 -500 9250 -300
rect 9450 -500 9600 -300
rect 9100 -600 9600 -500
rect 11600 -300 12100 -200
rect 11600 -500 11750 -300
rect 11950 -500 12100 -300
rect 11600 -600 12100 -500
rect 14100 -300 14600 -200
rect 14100 -500 14250 -300
rect 14450 -500 14600 -300
rect 14100 -600 14600 -500
rect 16600 -300 17100 -200
rect 16600 -500 16750 -300
rect 16950 -500 17100 -300
rect 16600 -600 17100 -500
rect 19100 -300 19600 -200
rect 19100 -500 19250 -300
rect 19450 -500 19600 -300
rect 19100 -600 19600 -500
rect 21600 -300 22100 -200
rect 21600 -500 21750 -300
rect 21950 -500 22100 -300
rect 21600 -600 22100 -500
rect 24100 -300 24600 -200
rect 24100 -500 24250 -300
rect 24450 -500 24600 -300
rect 24100 -600 24600 -500
rect 26600 -300 27100 -200
rect 26600 -500 26750 -300
rect 26950 -500 27100 -300
rect 26600 -600 27100 -500
rect 29100 -300 29600 -200
rect 29100 -500 29250 -300
rect 29450 -500 29600 -300
rect 29100 -600 29600 -500
rect 31600 -300 32000 -200
rect 31600 -500 31700 -300
rect 31900 -500 32000 -300
rect 31600 -600 32000 -500
rect 33200 -300 33600 -200
rect 33200 -500 33300 -300
rect 33500 -500 33600 -300
rect 33200 -600 33600 -500
<< nsubdiffcont >>
rect -800 2000 -600 2200
rect 1750 2000 1950 2200
rect 4250 2000 4450 2200
rect 6750 2000 6950 2200
rect 9250 2000 9450 2200
rect 11750 2000 11950 2200
rect 14250 2000 14450 2200
rect 16750 2000 16950 2200
rect 19250 2000 19450 2200
rect 21750 2000 21950 2200
rect 24250 2000 24450 2200
rect 26750 2000 26950 2200
rect 29250 2000 29450 2200
rect 31700 2000 31900 2200
rect 33300 2000 33500 2200
rect -800 -500 -600 -300
rect 1750 -500 1950 -300
rect 4250 -500 4450 -300
rect 6750 -500 6950 -300
rect 9250 -500 9450 -300
rect 11750 -500 11950 -300
rect 14250 -500 14450 -300
rect 16750 -500 16950 -300
rect 19250 -500 19450 -300
rect 21750 -500 21950 -300
rect 24250 -500 24450 -300
rect 26750 -500 26950 -300
rect 29250 -500 29450 -300
rect 31700 -500 31900 -300
rect 33300 -500 33500 -300
<< poly >>
rect 0 2300 1200 2335
rect 2500 2300 3700 2335
rect 5000 2300 6200 2335
rect 7500 2300 8700 2335
rect 10000 2300 11200 2335
rect 12500 2300 13700 2335
rect 15000 2300 16200 2335
rect 17500 2300 18700 2335
rect 20000 2300 21200 2335
rect 22500 2300 23700 2335
rect 25000 2300 26200 2335
rect 27500 2300 28700 2335
rect 30000 2300 31200 2335
rect 0 1800 1200 1900
rect 2500 1800 3700 1900
rect 5000 1800 6200 1900
rect 7500 1800 8700 1900
rect 10000 1800 11200 1900
rect 12500 1800 13700 1900
rect 15000 1800 16200 1900
rect 17500 1800 18700 1900
rect 20000 1800 21200 1900
rect 22500 1800 23700 1900
rect 25000 1800 26200 1900
rect 27500 1800 28700 1900
rect 30000 1800 31200 1900
rect 32000 1800 33200 1850
rect 0 1300 1200 1400
rect 2500 1300 3700 1400
rect 5000 1300 6200 1400
rect 7500 1300 8700 1400
rect 10000 1300 11200 1400
rect 12500 1300 13700 1400
rect 15000 1300 16200 1400
rect 17500 1300 18700 1400
rect 20000 1300 21200 1400
rect 22500 1300 23700 1400
rect 25000 1300 26200 1400
rect 27500 1300 28700 1400
rect 30000 1300 31200 1400
rect 32000 1300 33200 1400
rect -900 1200 -500 1300
rect -900 1000 -800 1200
rect -600 1000 -500 1200
rect -900 800 -500 1000
rect 0 800 1200 900
rect 2500 800 3700 900
rect 5000 800 6200 900
rect 7500 800 8700 900
rect 10000 800 11200 900
rect 12500 800 13700 900
rect 15000 800 16200 900
rect 17500 800 18700 900
rect 20000 800 21200 900
rect 22500 800 23700 900
rect 25000 800 26200 900
rect 27500 800 28700 900
rect 30000 800 31200 900
rect 32000 800 33200 900
rect -900 419 33200 800
rect -901 400 33200 419
rect 0 300 1200 400
rect 2500 300 3700 400
rect 5000 300 6200 400
rect 7500 300 8700 400
rect 10000 300 11200 400
rect 12500 300 13700 400
rect 15000 300 16200 400
rect 17500 300 18700 400
rect 20000 300 21200 400
rect 22500 300 23700 400
rect 25000 300 26200 400
rect 27500 300 28700 400
rect 30000 300 31200 400
rect 0 -200 1200 -100
rect 2500 -200 3700 -100
rect 5000 -200 6200 -100
rect 7500 -200 8700 -100
rect 10000 -200 11200 -100
rect 12500 -200 13700 -100
rect 15000 -200 16200 -100
rect 17500 -200 18700 -100
rect 20000 -200 21200 -100
rect 22500 -200 23700 -100
rect 25000 -200 26200 -100
rect 27500 -200 28700 -100
rect 30000 -200 31200 -100
rect 0 -635 1200 -600
rect 2500 -635 3700 -600
rect 5000 -635 6200 -600
rect 7500 -635 8700 -600
rect 10000 -635 11200 -600
rect 12500 -635 13700 -600
rect 15000 -635 16200 -600
rect 17500 -635 18700 -600
rect 20000 -635 21200 -600
rect 22500 -635 23700 -600
rect 25000 -635 26200 -600
rect 27500 -635 28700 -600
rect 30000 -635 31200 -600
<< polycont >>
rect -800 1000 -600 1200
<< locali >>
rect -900 2200 33600 2300
rect -900 2000 -800 2200
rect -600 2000 -300 2200
rect -100 2000 1300 2200
rect 1500 2000 1750 2200
rect 1950 2000 2200 2200
rect 2400 2000 3800 2200
rect 4000 2000 4250 2200
rect 4450 2000 4700 2200
rect 4900 2000 6300 2200
rect 6500 2000 6750 2200
rect 6950 2000 7200 2200
rect 7400 2000 8800 2200
rect 9000 2000 9250 2200
rect 9450 2000 9700 2200
rect 9900 2000 11300 2200
rect 11500 2000 11750 2200
rect 11950 2000 12200 2200
rect 12400 2000 13800 2200
rect 14000 2000 14250 2200
rect 14450 2000 14700 2200
rect 14900 2000 16300 2200
rect 16500 2000 16750 2200
rect 16950 2000 17200 2200
rect 17400 2000 18800 2200
rect 19000 2000 19250 2200
rect 19450 2000 19700 2200
rect 19900 2000 21300 2200
rect 21500 2000 21750 2200
rect 21950 2000 22200 2200
rect 22400 2000 23800 2200
rect 24000 2000 24250 2200
rect 24450 2000 24700 2200
rect 24900 2000 26300 2200
rect 26500 2000 26750 2200
rect 26950 2000 27200 2200
rect 27400 2000 28800 2200
rect 29000 2000 29250 2200
rect 29450 2000 29700 2200
rect 29900 2000 31300 2200
rect 31500 2000 31700 2200
rect 31900 2000 33300 2200
rect 33500 2000 33600 2200
rect -900 1900 33600 2000
rect -400 1700 0 1900
rect -400 1500 -300 1700
rect -100 1500 0 1700
rect -900 1200 -500 1300
rect -900 1000 -800 1200
rect -600 1000 -500 1200
rect -900 900 -500 1000
rect -400 1200 0 1500
rect -400 1000 -300 1200
rect -100 1000 0 1200
rect -400 800 0 1000
rect -900 419 0 800
rect -901 400 0 419
rect -400 200 0 400
rect -400 0 -300 200
rect -100 0 0 200
rect -400 -200 0 0
rect 400 -200 800 1900
rect 1200 1700 2000 1800
rect 1200 1500 1300 1700
rect 1500 1500 2000 1700
rect 1200 1200 2000 1500
rect 1200 1000 1300 1200
rect 1500 1000 2000 1200
rect 1200 900 2000 1000
rect 1600 800 2000 900
rect 2100 1700 2500 1800
rect 2100 1500 2200 1700
rect 2400 1500 2500 1700
rect 2100 1200 2500 1500
rect 2100 1000 2200 1200
rect 2400 1000 2500 1200
rect 2100 800 2500 1000
rect 1600 400 2500 800
rect 1200 200 2000 300
rect 1200 0 1300 200
rect 1500 0 1700 200
rect 1900 0 2000 200
rect 1200 -100 2000 0
rect 2100 200 2500 400
rect 2100 0 2200 200
rect 2400 0 2500 200
rect 2100 -100 2500 0
rect 2900 -200 3300 1900
rect 3700 1700 4500 1800
rect 3700 1500 3800 1700
rect 4000 1500 4500 1700
rect 3700 1200 4500 1500
rect 3700 1000 3800 1200
rect 4000 1000 4500 1200
rect 3700 900 4500 1000
rect 4100 800 4500 900
rect 4600 1700 5000 1800
rect 4600 1500 4700 1700
rect 4900 1500 5000 1700
rect 4600 1200 5000 1500
rect 4600 1000 4700 1200
rect 4900 1000 5000 1200
rect 4600 800 5000 1000
rect 4100 400 5000 800
rect 3700 200 4500 300
rect 3700 0 3800 200
rect 4000 0 4200 200
rect 4400 0 4500 200
rect 3700 -100 4500 0
rect 4600 200 5000 400
rect 4600 0 4700 200
rect 4900 0 5000 200
rect 4600 -100 5000 0
rect 5400 -200 5800 1900
rect 6200 1700 7000 1800
rect 6200 1500 6300 1700
rect 6500 1500 7000 1700
rect 6200 1200 7000 1500
rect 6200 1000 6300 1200
rect 6500 1000 7000 1200
rect 6200 900 7000 1000
rect 6600 800 7000 900
rect 7100 1700 7500 1800
rect 7100 1500 7200 1700
rect 7400 1500 7500 1700
rect 7100 1200 7500 1500
rect 7100 1000 7200 1200
rect 7400 1000 7500 1200
rect 7100 800 7500 1000
rect 6600 400 7500 800
rect 6200 200 7000 300
rect 6200 0 6300 200
rect 6500 0 6700 200
rect 6900 0 7000 200
rect 6200 -100 7000 0
rect 7100 200 7500 400
rect 7100 0 7200 200
rect 7400 0 7500 200
rect 7100 -100 7500 0
rect 7900 -200 8300 1900
rect 8700 1700 9500 1800
rect 8700 1500 8800 1700
rect 9000 1500 9500 1700
rect 8700 1200 9500 1500
rect 8700 1000 8800 1200
rect 9000 1000 9500 1200
rect 8700 900 9500 1000
rect 9100 800 9500 900
rect 9600 1700 10000 1800
rect 9600 1500 9700 1700
rect 9900 1500 10000 1700
rect 9600 1200 10000 1500
rect 9600 1000 9700 1200
rect 9900 1000 10000 1200
rect 9600 800 10000 1000
rect 9100 400 10000 800
rect 8700 200 9500 300
rect 8700 0 8800 200
rect 9000 0 9200 200
rect 9400 0 9500 200
rect 8700 -100 9500 0
rect 9600 200 10000 400
rect 9600 0 9700 200
rect 9900 0 10000 200
rect 9600 -100 10000 0
rect 10400 -200 10800 1900
rect 11200 1700 12000 1800
rect 11200 1500 11300 1700
rect 11500 1500 12000 1700
rect 11200 1200 12000 1500
rect 11200 1000 11300 1200
rect 11500 1000 12000 1200
rect 11200 900 12000 1000
rect 11600 800 12000 900
rect 12100 1700 12500 1800
rect 12100 1500 12200 1700
rect 12400 1500 12500 1700
rect 12100 1200 12500 1500
rect 12100 1000 12200 1200
rect 12400 1000 12500 1200
rect 12100 800 12500 1000
rect 11600 400 12500 800
rect 11200 200 12000 300
rect 11200 0 11300 200
rect 11500 0 11700 200
rect 11900 0 12000 200
rect 11200 -100 12000 0
rect 12100 200 12500 400
rect 12100 0 12200 200
rect 12400 0 12500 200
rect 12100 -100 12500 0
rect 12900 -200 13300 1900
rect 13700 1700 14500 1800
rect 13700 1500 13800 1700
rect 14000 1500 14500 1700
rect 13700 1200 14500 1500
rect 13700 1000 13800 1200
rect 14000 1000 14500 1200
rect 13700 900 14500 1000
rect 14100 800 14500 900
rect 14600 1700 15000 1800
rect 14600 1500 14700 1700
rect 14900 1500 15000 1700
rect 14600 1200 15000 1500
rect 14600 1000 14700 1200
rect 14900 1000 15000 1200
rect 14600 800 15000 1000
rect 14100 400 15000 800
rect 13700 200 14500 300
rect 13700 0 13800 200
rect 14000 0 14200 200
rect 14400 0 14500 200
rect 13700 -100 14500 0
rect 14600 200 15000 400
rect 14600 0 14700 200
rect 14900 0 15000 200
rect 14600 -100 15000 0
rect 15400 -200 15800 1900
rect 16200 1700 17000 1800
rect 16200 1500 16300 1700
rect 16500 1500 17000 1700
rect 16200 1200 17000 1500
rect 16200 1000 16300 1200
rect 16500 1000 17000 1200
rect 16200 900 17000 1000
rect 16600 800 17000 900
rect 17100 1700 17500 1800
rect 17100 1500 17200 1700
rect 17400 1500 17500 1700
rect 17100 1200 17500 1500
rect 17100 1000 17200 1200
rect 17400 1000 17500 1200
rect 17100 800 17500 1000
rect 16600 400 17500 800
rect 16200 200 17000 300
rect 16200 0 16300 200
rect 16500 0 16700 200
rect 16900 0 17000 200
rect 16200 -100 17000 0
rect 17100 200 17500 400
rect 17100 0 17200 200
rect 17400 0 17500 200
rect 17100 -100 17500 0
rect 17900 -200 18300 1900
rect 18700 1700 19500 1800
rect 18700 1500 18800 1700
rect 19000 1500 19500 1700
rect 18700 1200 19500 1500
rect 18700 1000 18800 1200
rect 19000 1000 19500 1200
rect 18700 900 19500 1000
rect 19100 800 19500 900
rect 19600 1700 20000 1800
rect 19600 1500 19700 1700
rect 19900 1500 20000 1700
rect 19600 1200 20000 1500
rect 19600 1000 19700 1200
rect 19900 1000 20000 1200
rect 19600 800 20000 1000
rect 19100 400 20000 800
rect 18700 200 19500 300
rect 18700 0 18800 200
rect 19000 0 19200 200
rect 19400 0 19500 200
rect 18700 -100 19500 0
rect 19600 200 20000 400
rect 19600 0 19700 200
rect 19900 0 20000 200
rect 19600 -100 20000 0
rect 20400 -200 20800 1900
rect 21200 1700 22000 1800
rect 21200 1500 21300 1700
rect 21500 1500 22000 1700
rect 21200 1200 22000 1500
rect 21200 1000 21300 1200
rect 21500 1000 22000 1200
rect 21200 900 22000 1000
rect 21600 800 22000 900
rect 22100 1700 22500 1800
rect 22100 1500 22200 1700
rect 22400 1500 22500 1700
rect 22100 1200 22500 1500
rect 22100 1000 22200 1200
rect 22400 1000 22500 1200
rect 22100 800 22500 1000
rect 21600 400 22500 800
rect 21200 200 22000 300
rect 21200 0 21300 200
rect 21500 0 21700 200
rect 21900 0 22000 200
rect 21200 -100 22000 0
rect 22100 200 22500 400
rect 22100 0 22200 200
rect 22400 0 22500 200
rect 22100 -100 22500 0
rect 22900 -200 23300 1900
rect 23700 1700 24500 1800
rect 23700 1500 23800 1700
rect 24000 1500 24500 1700
rect 23700 1200 24500 1500
rect 23700 1000 23800 1200
rect 24000 1000 24500 1200
rect 23700 900 24500 1000
rect 24100 800 24500 900
rect 24600 1700 25000 1800
rect 24600 1500 24700 1700
rect 24900 1500 25000 1700
rect 24600 1200 25000 1500
rect 24600 1000 24700 1200
rect 24900 1000 25000 1200
rect 24600 800 25000 1000
rect 24100 400 25000 800
rect 23700 200 24500 300
rect 23700 0 23800 200
rect 24000 0 24200 200
rect 24400 0 24500 200
rect 23700 -100 24500 0
rect 24600 200 25000 400
rect 24600 0 24700 200
rect 24900 0 25000 200
rect 24600 -100 25000 0
rect 25400 -200 25800 1900
rect 26200 1700 27000 1800
rect 26200 1500 26300 1700
rect 26500 1500 27000 1700
rect 26200 1200 27000 1500
rect 26200 1000 26300 1200
rect 26500 1000 27000 1200
rect 26200 900 27000 1000
rect 26600 800 27000 900
rect 27100 1700 27500 1800
rect 27100 1500 27200 1700
rect 27400 1500 27500 1700
rect 27100 1200 27500 1500
rect 27100 1000 27200 1200
rect 27400 1000 27500 1200
rect 27100 800 27500 1000
rect 26600 400 27500 800
rect 26200 200 27000 300
rect 26200 0 26300 200
rect 26500 0 26700 200
rect 26900 0 27000 200
rect 26200 -100 27000 0
rect 27100 200 27500 400
rect 27100 0 27200 200
rect 27400 0 27500 200
rect 27100 -100 27500 0
rect 27900 -200 28300 1900
rect 28700 1700 29500 1800
rect 28700 1500 28800 1700
rect 29000 1500 29500 1700
rect 28700 1200 29500 1500
rect 28700 1000 28800 1200
rect 29000 1000 29500 1200
rect 28700 900 29500 1000
rect 29100 800 29500 900
rect 29600 1700 30000 1800
rect 29600 1500 29700 1700
rect 29900 1500 30000 1700
rect 29600 1200 30000 1500
rect 29600 1000 29700 1200
rect 29900 1000 30000 1200
rect 29600 800 30000 1000
rect 29100 400 30000 800
rect 28700 200 29500 300
rect 28700 0 28800 200
rect 29000 0 29200 200
rect 29400 0 29500 200
rect 28700 -100 29500 0
rect 29600 200 30000 400
rect 29600 0 29700 200
rect 29900 0 30000 200
rect 29600 -100 30000 0
rect 30400 -200 30800 1900
rect 31200 1700 32000 1800
rect 31200 1500 31300 1700
rect 31500 1500 31700 1700
rect 31900 1500 32000 1700
rect 31200 1200 32000 1500
rect 31200 1000 31300 1200
rect 31500 1000 31700 1200
rect 31900 1000 32000 1200
rect 31200 900 32000 1000
rect 33200 1700 33600 1800
rect 33200 1500 33300 1700
rect 33500 1500 33600 1700
rect 33200 1200 33600 1500
rect 33200 1000 33300 1200
rect 33500 1000 33600 1200
rect 33200 400 33600 1000
rect 31200 200 32000 300
rect 31200 0 31300 200
rect 31500 0 31700 200
rect 31900 0 32000 200
rect 31200 -100 32000 0
rect -900 -300 33600 -200
rect -900 -500 -800 -300
rect -600 -500 -300 -300
rect -100 -500 1300 -300
rect 1500 -500 1750 -300
rect 1950 -500 2200 -300
rect 2400 -500 3800 -300
rect 4000 -500 4250 -300
rect 4450 -500 4700 -300
rect 4900 -500 6300 -300
rect 6500 -500 6750 -300
rect 6950 -500 7200 -300
rect 7400 -500 8800 -300
rect 9000 -500 9250 -300
rect 9450 -500 9700 -300
rect 9900 -500 11300 -300
rect 11500 -500 11750 -300
rect 11950 -500 12200 -300
rect 12400 -500 13800 -300
rect 14000 -500 14250 -300
rect 14450 -500 14700 -300
rect 14900 -500 16300 -300
rect 16500 -500 16750 -300
rect 16950 -500 17200 -300
rect 17400 -500 18800 -300
rect 19000 -500 19250 -300
rect 19450 -500 19700 -300
rect 19900 -500 21300 -300
rect 21500 -500 21750 -300
rect 21950 -500 22200 -300
rect 22400 -500 23800 -300
rect 24000 -500 24250 -300
rect 24450 -500 24700 -300
rect 24900 -500 26300 -300
rect 26500 -500 26750 -300
rect 26950 -500 27200 -300
rect 27400 -500 28800 -300
rect 29000 -500 29250 -300
rect 29450 -500 29700 -300
rect 29900 -500 31300 -300
rect 31500 -500 31700 -300
rect 31900 -500 33300 -300
rect 33500 -500 33600 -300
rect -900 -600 33600 -500
<< viali >>
rect 1700 0 1900 200
rect 4200 0 4400 200
rect 6700 0 6900 200
rect 9200 0 9400 200
rect 11700 0 11900 200
rect 14200 0 14400 200
rect 16700 0 16900 200
rect 19200 0 19400 200
rect 21700 0 21900 200
rect 24200 0 24400 200
rect 26700 0 26900 200
rect 29200 0 29400 200
rect 31700 0 31900 200
<< metal1 >>
rect 1600 200 2000 300
rect 1600 0 1700 200
rect 1900 0 2000 200
rect 1600 -600 2000 0
rect 4100 200 4500 300
rect 4100 0 4200 200
rect 4400 0 4500 200
rect 4100 -600 4500 0
rect 6600 200 7000 300
rect 6600 0 6700 200
rect 6900 0 7000 200
rect 6600 -600 7000 0
rect 9100 200 9500 300
rect 9100 0 9200 200
rect 9400 0 9500 200
rect 9100 -600 9500 0
rect 11600 200 12000 300
rect 11600 0 11700 200
rect 11900 0 12000 200
rect 11600 -600 12000 0
rect 14100 200 14500 300
rect 14100 0 14200 200
rect 14400 0 14500 200
rect 14100 -600 14500 0
rect 16600 200 17000 300
rect 16600 0 16700 200
rect 16900 0 17000 200
rect 16600 -600 17000 0
rect 19100 200 19500 300
rect 19100 0 19200 200
rect 19400 0 19500 200
rect 19100 -600 19500 0
rect 21600 200 22000 300
rect 21600 0 21700 200
rect 21900 0 22000 200
rect 21600 -600 22000 0
rect 24100 200 24500 300
rect 24100 0 24200 200
rect 24400 0 24500 200
rect 24100 -600 24500 0
rect 26600 200 27000 300
rect 26600 0 26700 200
rect 26900 0 27000 200
rect 26600 -600 27000 0
rect 29100 200 29500 300
rect 29100 0 29200 200
rect 29400 0 29500 200
rect 29100 -600 29500 0
rect 31600 200 32000 300
rect 31600 0 31700 200
rect 31900 0 32000 200
rect 31600 -600 32000 0
rect -900 -1000 32000 -600
<< labels >>
rlabel locali -900 900 -900 1300 7 VGATE
port 2 w
rlabel nwell -900 400 -900 800 7 VP
port 3 w
rlabel metal1 -900 -1000 -900 -600 7 VN
port 4 w
rlabel locali 33600 400 33600 800 3 IOUT
port 5 e
<< end >>
